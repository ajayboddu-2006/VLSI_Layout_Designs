magic
tech sky130A
timestamp 1737365683
<< nwell >>
rect -361 493 -63 494
rect -361 492 882 493
rect -361 247 971 492
<< nmos >>
rect -255 27 -240 86
rect -128 27 -113 86
rect 0 27 15 88
rect 58 27 73 88
rect 118 27 133 88
rect 178 27 193 88
rect 238 27 253 88
rect 298 27 313 88
rect 358 27 373 88
rect 418 27 433 88
rect 478 27 493 88
rect 538 27 553 88
rect 598 27 613 88
rect 658 27 673 88
rect 804 26 819 87
<< pmos >>
rect -255 267 -240 327
rect -128 267 -113 327
rect 0 267 15 328
rect 58 267 73 328
rect 118 267 133 328
rect 178 267 193 328
rect 238 267 253 328
rect 298 267 313 328
rect 358 267 373 328
rect 418 267 433 328
rect 478 267 493 328
rect 538 267 553 328
rect 598 267 613 328
rect 658 267 673 328
rect 804 267 819 328
<< ndiff >>
rect -298 78 -255 86
rect -298 38 -284 78
rect -263 38 -255 78
rect -298 27 -255 38
rect -240 78 -198 86
rect -240 38 -226 78
rect -205 38 -198 78
rect -240 27 -198 38
rect -171 79 -128 86
rect -171 39 -159 79
rect -138 39 -128 79
rect -171 27 -128 39
rect -113 78 -70 86
rect -113 38 -100 78
rect -79 38 -70 78
rect -113 27 -70 38
rect -43 77 0 88
rect -43 37 -32 77
rect -11 37 0 77
rect -43 27 0 37
rect 15 27 58 88
rect 73 27 118 88
rect 133 78 178 88
rect 133 38 147 78
rect 168 38 178 78
rect 133 27 178 38
rect 193 27 238 88
rect 253 27 298 88
rect 313 78 358 88
rect 313 38 325 78
rect 346 38 358 78
rect 313 27 358 38
rect 373 27 418 88
rect 433 27 478 88
rect 493 78 538 88
rect 493 38 506 78
rect 527 38 538 78
rect 493 27 538 38
rect 553 27 598 88
rect 613 27 658 88
rect 673 79 718 88
rect 673 39 686 79
rect 707 39 718 79
rect 673 27 718 39
rect 760 81 804 87
rect 760 41 774 81
rect 795 41 804 81
rect 760 26 804 41
rect 819 77 863 87
rect 819 37 833 77
rect 854 37 863 77
rect 819 26 863 37
<< pdiff >>
rect -297 320 -255 327
rect -297 280 -285 320
rect -265 280 -255 320
rect -297 267 -255 280
rect -240 320 -197 327
rect -240 280 -227 320
rect -207 280 -197 320
rect -240 267 -197 280
rect -170 318 -128 327
rect -170 278 -160 318
rect -140 278 -128 318
rect -170 267 -128 278
rect -113 318 -70 327
rect -113 278 -100 318
rect -80 278 -70 318
rect -113 267 -70 278
rect -43 318 0 328
rect -43 278 -32 318
rect -12 278 0 318
rect -43 267 0 278
rect 15 319 58 328
rect 15 279 28 319
rect 48 279 58 319
rect 15 267 58 279
rect 73 319 118 328
rect 73 279 88 319
rect 108 279 118 319
rect 73 267 118 279
rect 133 320 178 328
rect 133 280 146 320
rect 166 280 178 320
rect 133 267 178 280
rect 193 319 238 328
rect 193 279 205 319
rect 225 279 238 319
rect 193 267 238 279
rect 253 319 298 328
rect 253 279 267 319
rect 287 279 298 319
rect 253 267 298 279
rect 313 319 358 328
rect 313 279 328 319
rect 348 279 358 319
rect 313 267 358 279
rect 373 318 418 328
rect 373 278 388 318
rect 408 278 418 318
rect 373 267 418 278
rect 433 319 478 328
rect 433 279 447 319
rect 467 279 478 319
rect 433 267 478 279
rect 493 318 538 328
rect 493 278 507 318
rect 527 278 538 318
rect 493 267 538 278
rect 553 318 598 328
rect 553 278 568 318
rect 588 278 598 318
rect 553 267 598 278
rect 613 317 658 328
rect 613 277 626 317
rect 646 277 658 317
rect 613 267 658 277
rect 673 317 718 328
rect 673 277 685 317
rect 705 277 718 317
rect 673 267 718 277
rect 759 318 804 328
rect 759 278 774 318
rect 794 278 804 318
rect 759 267 804 278
rect 819 320 864 328
rect 819 280 832 320
rect 852 280 864 320
rect 819 267 864 280
<< ndiffc >>
rect -284 38 -263 78
rect -226 38 -205 78
rect -159 39 -138 79
rect -100 38 -79 78
rect -32 37 -11 77
rect 147 38 168 78
rect 325 38 346 78
rect 506 38 527 78
rect 686 39 707 79
rect 774 41 795 81
rect 833 37 854 77
<< pdiffc >>
rect -285 280 -265 320
rect -227 280 -207 320
rect -160 278 -140 318
rect -100 278 -80 318
rect -32 278 -12 318
rect 28 279 48 319
rect 88 279 108 319
rect 146 280 166 320
rect 205 279 225 319
rect 267 279 287 319
rect 328 279 348 319
rect 388 278 408 318
rect 447 279 467 319
rect 507 278 527 318
rect 568 278 588 318
rect 626 277 646 317
rect 685 277 705 317
rect 774 278 794 318
rect 832 280 852 320
<< psubdiff >>
rect -355 -44 951 -36
rect -355 -47 128 -44
rect -355 -70 9 -47
rect 33 -50 128 -47
rect 33 -70 75 -50
rect -355 -73 75 -70
rect 99 -67 128 -50
rect 152 -46 387 -44
rect 152 -67 197 -46
rect 99 -69 197 -67
rect 221 -47 387 -46
rect 221 -69 262 -47
rect 99 -70 262 -69
rect 286 -67 387 -47
rect 411 -46 511 -44
rect 411 -67 448 -46
rect 286 -69 448 -67
rect 472 -67 511 -46
rect 535 -48 951 -44
rect 535 -67 580 -48
rect 472 -69 580 -67
rect 286 -70 580 -69
rect 99 -71 580 -70
rect 604 -71 639 -48
rect 663 -71 951 -48
rect 99 -73 951 -71
rect -355 -84 951 -73
<< nsubdiff >>
rect -342 449 953 460
rect -342 447 148 449
rect -342 424 20 447
rect 44 426 148 447
rect 172 448 335 449
rect 172 447 271 448
rect 172 426 210 447
rect 44 424 210 426
rect 234 425 271 447
rect 295 426 335 448
rect 359 447 462 449
rect 359 426 396 447
rect 295 425 396 426
rect 234 424 396 425
rect 420 426 462 447
rect 486 447 661 449
rect 486 426 523 447
rect 420 424 523 426
rect 547 424 597 447
rect 621 426 661 447
rect 685 426 953 449
rect 621 424 953 426
rect -342 412 953 424
<< psubdiffcont >>
rect 9 -70 33 -47
rect 75 -73 99 -50
rect 128 -67 152 -44
rect 197 -69 221 -46
rect 262 -70 286 -47
rect 387 -67 411 -44
rect 448 -69 472 -46
rect 511 -67 535 -44
rect 580 -71 604 -48
rect 639 -71 663 -48
<< nsubdiffcont >>
rect 20 424 44 447
rect 148 426 172 449
rect 210 424 234 447
rect 271 425 295 448
rect 335 426 359 449
rect 396 424 420 447
rect 462 426 486 449
rect 523 424 547 447
rect 597 424 621 447
rect 661 426 685 449
<< poly >>
rect -255 327 -240 370
rect -128 327 -113 371
rect 0 328 15 369
rect 58 328 73 369
rect 118 328 133 369
rect 178 328 193 369
rect 238 328 253 369
rect 298 328 313 369
rect 358 328 373 369
rect 418 328 433 369
rect 478 328 493 369
rect 538 328 553 369
rect 598 328 613 369
rect 658 328 673 369
rect 804 328 819 369
rect -255 189 -240 267
rect -272 166 -240 189
rect -128 175 -113 267
rect -255 86 -240 166
rect -152 152 -113 175
rect -128 86 -113 152
rect 0 88 15 267
rect 58 189 73 267
rect 118 247 133 267
rect 178 247 193 267
rect 108 239 140 247
rect 108 222 116 239
rect 133 222 140 239
rect 108 214 140 222
rect 174 239 206 247
rect 174 222 181 239
rect 198 222 206 239
rect 174 214 206 222
rect 48 181 81 189
rect 48 164 56 181
rect 73 164 81 181
rect 48 156 81 164
rect 58 88 73 156
rect 118 88 133 214
rect 178 88 193 214
rect 238 88 253 267
rect 298 88 313 267
rect 358 88 373 267
rect 418 187 433 267
rect 409 179 441 187
rect 409 162 419 179
rect 436 162 441 179
rect 409 154 441 162
rect 418 88 433 154
rect 478 88 493 267
rect 538 88 553 267
rect 598 88 613 267
rect 658 88 673 267
rect 750 130 783 138
rect 804 130 819 267
rect 750 113 758 130
rect 775 113 819 130
rect 750 105 783 113
rect 804 87 819 113
rect -255 -4 -240 27
rect -128 -4 -113 27
rect 0 -4 15 27
rect 58 -4 73 27
rect 118 -4 133 27
rect 178 -4 193 27
rect 238 -4 253 27
rect 298 -4 313 27
rect 358 -4 373 27
rect 418 -4 433 27
rect 478 -4 493 27
rect 538 -4 553 27
rect 598 -4 613 27
rect 658 -4 673 27
rect 804 -2 819 26
<< polycont >>
rect 116 222 133 239
rect 181 222 198 239
rect 56 164 73 181
rect 419 162 436 179
rect 758 113 775 130
<< locali >>
rect -361 450 971 460
rect -361 449 710 450
rect -361 447 148 449
rect -361 445 -164 447
rect -361 422 -337 445
rect -313 422 -286 445
rect -262 422 -229 445
rect -205 424 -164 445
rect -140 424 -103 447
rect -79 445 20 447
rect -79 424 -46 445
rect -205 422 -46 424
rect -22 424 20 445
rect 44 446 148 447
rect 44 424 87 446
rect -22 423 87 424
rect 111 426 148 446
rect 172 448 335 449
rect 172 447 271 448
rect 172 426 210 447
rect 111 424 210 426
rect 234 425 271 447
rect 295 426 335 448
rect 359 447 462 449
rect 359 426 396 447
rect 295 425 396 426
rect 234 424 396 425
rect 420 426 462 447
rect 486 447 661 449
rect 486 426 523 447
rect 420 424 523 426
rect 547 424 597 447
rect 621 426 661 447
rect 685 427 710 449
rect 734 448 971 450
rect 734 427 765 448
rect 685 426 765 427
rect 621 425 765 426
rect 789 425 819 448
rect 843 447 971 448
rect 843 425 888 447
rect 621 424 888 425
rect 912 424 971 447
rect 111 423 971 424
rect -22 422 971 423
rect -361 412 971 422
rect -286 327 -264 412
rect -159 327 -137 412
rect -43 328 -22 412
rect 88 328 109 412
rect 204 345 467 366
rect 204 328 225 345
rect 327 328 348 345
rect 446 328 467 345
rect 764 328 792 412
rect -297 320 -257 327
rect -297 280 -285 320
rect -265 280 -257 320
rect -297 267 -257 280
rect -238 320 -197 327
rect -238 280 -227 320
rect -207 280 -197 320
rect -238 267 -197 280
rect -170 318 -130 327
rect -170 278 -160 318
rect -140 278 -130 318
rect -170 267 -130 278
rect -111 318 -70 327
rect -111 278 -100 318
rect -80 278 -70 318
rect -111 267 -70 278
rect -43 318 -2 328
rect -43 278 -32 318
rect -12 278 -2 318
rect -43 267 -2 278
rect 16 319 57 328
rect 16 279 28 319
rect 48 279 57 319
rect 16 267 57 279
rect 74 319 117 328
rect 74 279 88 319
rect 108 279 117 319
rect 74 267 117 279
rect 134 320 177 328
rect 134 280 146 320
rect 166 280 177 320
rect 134 267 177 280
rect 194 319 237 328
rect 194 279 205 319
rect 225 279 237 319
rect 194 267 237 279
rect 254 319 297 328
rect 254 279 267 319
rect 287 279 297 319
rect 254 267 297 279
rect 314 319 357 328
rect 314 279 328 319
rect 348 279 357 319
rect 314 267 357 279
rect 374 318 417 328
rect 374 278 388 318
rect 408 278 417 318
rect 374 267 417 278
rect 434 319 477 328
rect 434 279 447 319
rect 467 279 477 319
rect 434 267 477 279
rect 494 318 537 328
rect 494 278 507 318
rect 527 278 537 318
rect 494 267 537 278
rect 554 318 597 328
rect 554 278 568 318
rect 588 278 597 318
rect 554 267 597 278
rect 614 317 657 328
rect 614 277 626 317
rect 646 277 657 317
rect 614 267 657 277
rect 674 317 718 328
rect 674 277 685 317
rect 705 277 718 317
rect 674 267 718 277
rect 759 318 803 328
rect 759 278 774 318
rect 794 278 803 318
rect 759 267 803 278
rect 820 320 864 328
rect 820 280 832 320
rect 852 280 864 320
rect 820 267 864 280
rect -226 240 -205 267
rect -182 240 -147 246
rect -226 223 -174 240
rect -155 223 -147 240
rect -226 86 -205 223
rect -182 215 -147 223
rect -100 180 -79 267
rect -62 239 -27 246
rect 108 239 140 247
rect 174 239 206 247
rect -62 222 -55 239
rect -36 222 116 239
rect 133 222 181 239
rect 198 222 206 239
rect -62 215 -27 222
rect 108 214 140 222
rect 174 214 206 222
rect 48 181 81 189
rect 48 180 56 181
rect -100 164 56 180
rect 73 180 81 181
rect 409 180 441 187
rect 73 179 441 180
rect 73 164 419 179
rect -100 163 419 164
rect -100 86 -79 163
rect 48 156 81 163
rect 409 162 419 163
rect 436 162 441 179
rect 409 154 441 162
rect 567 134 585 267
rect 689 134 707 267
rect 836 188 863 267
rect 836 165 882 188
rect 143 128 172 134
rect 143 111 150 128
rect 167 111 172 128
rect 143 105 172 111
rect 503 127 532 134
rect 503 110 509 127
rect 526 110 532 127
rect 503 105 532 110
rect 560 128 592 134
rect 560 111 568 128
rect 585 111 592 128
rect 560 105 592 111
rect 684 128 713 134
rect 750 130 783 138
rect 750 128 758 130
rect 684 111 691 128
rect 708 113 758 128
rect 775 113 783 130
rect 708 111 783 113
rect 684 105 713 111
rect 750 105 783 111
rect 150 88 167 105
rect 507 88 525 105
rect -298 78 -256 86
rect -298 38 -284 78
rect -263 38 -256 78
rect -298 27 -256 38
rect -239 78 -198 86
rect -239 38 -226 78
rect -205 38 -198 78
rect -239 27 -198 38
rect -171 79 -129 86
rect -171 39 -159 79
rect -138 39 -129 79
rect -171 27 -129 39
rect -112 78 -70 86
rect -112 38 -100 78
rect -79 38 -70 78
rect -112 27 -70 38
rect -43 77 -2 88
rect -43 37 -32 77
rect -11 37 -2 77
rect -43 27 -2 37
rect 135 78 176 88
rect 135 38 147 78
rect 168 38 176 78
rect 135 27 176 38
rect 315 78 356 88
rect 315 38 325 78
rect 346 38 356 78
rect 315 27 356 38
rect 495 78 536 88
rect 495 38 506 78
rect 527 38 536 78
rect 495 27 536 38
rect 675 79 718 88
rect 836 87 863 165
rect 675 39 686 79
rect 707 39 718 79
rect 675 27 718 39
rect -293 -36 -271 27
rect -161 -36 -139 27
rect -43 -36 -26 27
rect 325 -36 346 27
rect 697 -36 718 27
rect 760 81 803 87
rect 760 41 774 81
rect 795 41 803 81
rect 760 26 803 41
rect 820 77 863 87
rect 820 37 833 77
rect 854 37 863 77
rect 820 26 863 37
rect 767 -36 795 26
rect -355 -42 951 -36
rect -355 -44 -48 -42
rect -355 -47 -295 -44
rect -355 -70 -342 -47
rect -318 -67 -295 -47
rect -271 -67 -234 -44
rect -210 -47 -48 -44
rect -210 -50 -100 -47
rect -210 -67 -160 -50
rect -318 -70 -160 -67
rect -355 -73 -160 -70
rect -136 -70 -100 -50
rect -76 -65 -48 -47
rect -24 -44 324 -42
rect -24 -47 128 -44
rect -24 -65 9 -47
rect -76 -70 9 -65
rect 33 -50 128 -47
rect 33 -70 75 -50
rect -136 -73 75 -70
rect 99 -67 128 -50
rect 152 -46 324 -44
rect 152 -67 197 -46
rect 99 -69 197 -67
rect 221 -47 324 -46
rect 221 -69 262 -47
rect 99 -70 262 -69
rect 286 -65 324 -47
rect 348 -44 951 -42
rect 348 -65 387 -44
rect 286 -67 387 -65
rect 411 -46 511 -44
rect 411 -67 448 -46
rect 286 -69 448 -67
rect 472 -67 511 -46
rect 535 -47 951 -44
rect 535 -48 694 -47
rect 535 -67 580 -48
rect 472 -69 580 -67
rect 286 -70 580 -69
rect 99 -71 580 -70
rect 604 -71 639 -48
rect 663 -70 694 -48
rect 718 -48 838 -47
rect 718 -70 767 -48
rect 663 -71 767 -70
rect 791 -70 838 -48
rect 862 -70 897 -47
rect 921 -70 951 -47
rect 791 -71 951 -70
rect 99 -73 951 -71
rect -355 -84 951 -73
<< viali >>
rect -337 422 -313 445
rect -286 422 -262 445
rect -229 422 -205 445
rect -164 424 -140 447
rect -103 424 -79 447
rect -46 422 -22 445
rect 87 423 111 446
rect 710 427 734 450
rect 765 425 789 448
rect 819 425 843 448
rect 888 424 912 447
rect 28 279 48 319
rect 146 280 166 320
rect 267 279 287 319
rect 388 278 408 318
rect 507 278 527 318
rect 626 277 646 317
rect -174 223 -155 240
rect -55 222 -36 239
rect 150 111 167 128
rect 509 110 526 127
rect 568 111 585 128
rect 691 111 708 128
rect -342 -70 -318 -47
rect -295 -67 -271 -44
rect -234 -67 -210 -44
rect -160 -73 -136 -50
rect -100 -70 -76 -47
rect -48 -65 -24 -42
rect 324 -65 348 -42
rect 694 -70 718 -47
rect 767 -71 791 -48
rect 838 -70 862 -47
rect 897 -70 921 -47
<< metal1 >>
rect -361 450 971 460
rect -361 447 710 450
rect -361 445 -164 447
rect -361 422 -337 445
rect -313 422 -286 445
rect -262 422 -229 445
rect -205 424 -164 445
rect -140 424 -103 447
rect -79 446 710 447
rect -79 445 87 446
rect -79 424 -46 445
rect -205 422 -46 424
rect -22 423 87 445
rect 111 427 710 446
rect 734 448 971 450
rect 734 427 765 448
rect 111 425 765 427
rect 789 425 819 448
rect 843 447 971 448
rect 843 425 888 447
rect 111 424 888 425
rect 912 424 971 447
rect 111 423 971 424
rect -22 422 971 423
rect -361 412 971 422
rect 16 319 57 328
rect 16 279 28 319
rect 48 307 57 319
rect 134 320 177 328
rect 134 307 146 320
rect 48 289 146 307
rect 48 279 57 289
rect 16 267 57 279
rect 134 280 146 289
rect 166 307 177 320
rect 254 319 297 328
rect 254 307 267 319
rect 166 289 267 307
rect 166 280 177 289
rect 134 267 177 280
rect 254 279 267 289
rect 287 279 297 319
rect 254 267 297 279
rect 374 318 417 328
rect 374 278 388 318
rect 408 308 417 318
rect 494 318 537 328
rect 494 308 507 318
rect 408 290 507 308
rect 408 278 417 290
rect 374 267 417 278
rect 494 278 507 290
rect 527 308 537 318
rect 614 317 657 328
rect 614 308 626 317
rect 527 290 626 308
rect 527 278 537 290
rect 494 267 537 278
rect 614 277 626 290
rect 646 277 657 317
rect 614 267 657 277
rect -182 240 -147 246
rect -182 223 -174 240
rect -155 239 -147 240
rect -62 239 -27 246
rect -155 223 -55 239
rect -182 215 -147 223
rect -62 222 -55 223
rect -36 222 -27 239
rect -62 215 -27 222
rect 143 128 172 134
rect 143 111 150 128
rect 167 126 172 128
rect 503 127 532 134
rect 503 126 509 127
rect 167 112 509 126
rect 167 111 172 112
rect 143 105 172 111
rect 503 110 509 112
rect 526 126 532 127
rect 560 128 592 134
rect 560 126 568 128
rect 526 112 568 126
rect 526 110 532 112
rect 503 105 532 110
rect 560 111 568 112
rect 585 126 592 128
rect 684 128 713 134
rect 684 126 691 128
rect 585 112 691 126
rect 585 111 592 112
rect 560 105 592 111
rect 684 111 691 112
rect 708 111 713 128
rect 684 105 713 111
rect -355 -42 951 -36
rect -355 -44 -48 -42
rect -355 -47 -295 -44
rect -355 -70 -342 -47
rect -318 -67 -295 -47
rect -271 -67 -234 -44
rect -210 -47 -48 -44
rect -210 -50 -100 -47
rect -210 -67 -160 -50
rect -318 -70 -160 -67
rect -355 -73 -160 -70
rect -136 -70 -100 -50
rect -76 -65 -48 -47
rect -24 -65 324 -42
rect 348 -47 951 -42
rect 348 -65 694 -47
rect -76 -70 694 -65
rect 718 -48 838 -47
rect 718 -70 767 -48
rect -136 -71 767 -70
rect 791 -70 838 -48
rect 862 -70 897 -47
rect 921 -70 951 -47
rect 791 -71 951 -70
rect -136 -73 951 -71
rect -355 -84 951 -73
<< labels >>
flabel metal1 s -363 409 -313 461 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel metal1 s -350 -84 -300 -32 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel poly s -11 -6 24 23 0 FreeSans 80 0 0 0 I0
port 2 nsew
flabel poly s 288 -7 323 22 0 FreeSans 80 0 0 0 I1
port 3 nsew
flabel poly s 351 -7 386 22 0 FreeSans 80 0 0 0 I2
port 4 nsew
flabel poly s 651 -9 686 20 0 FreeSans 80 0 0 0 I3
port 5 nsew
flabel poly s -275 162 -240 191 0 FreeSans 80 0 0 0 S0
port 6 nsew
flabel poly s 471 -7 506 22 0 FreeSans 80 0 0 0 S0
flabel poly s 535 -7 570 22 0 FreeSans 80 0 0 0 S0
flabel poly s -157 148 -122 177 0 FreeSans 80 0 0 0 S1
port 7 nsew
flabel poly s 232 -8 267 21 0 FreeSans 80 0 0 0 S1
flabel poly s 591 -10 626 19 0 FreeSans 80 0 0 0 S1
flabel locali s 859 162 894 191 0 FreeSans 80 0 0 0 OUT
port 8 nsew
<< end >>
