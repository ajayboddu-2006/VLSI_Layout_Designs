magic
tech sky130A
timestamp 1737724314
<< nwell >>
rect -638 -886 1437 -678
rect -509 -1438 1457 -1230
<< nmos >>
rect -574 -1132 -557 -1067
rect -437 -1132 -420 -1067
rect -289 -1132 -272 -1067
rect -220 -1132 -203 -1067
rect -149 -1132 -132 -1067
rect -4 -1132 13 -1067
rect 163 -1132 180 -1067
rect 232 -1132 249 -1067
rect 303 -1132 320 -1067
rect 448 -1132 465 -1067
rect 618 -1132 635 -1067
rect 687 -1132 704 -1067
rect 758 -1132 775 -1067
rect 903 -1132 920 -1067
rect 1068 -1132 1085 -1067
rect 1137 -1132 1154 -1067
rect 1208 -1132 1225 -1067
rect 1353 -1132 1370 -1067
rect -445 -1684 -428 -1619
rect -293 -1684 -276 -1619
rect -224 -1684 -207 -1619
rect -153 -1684 -136 -1619
rect -8 -1684 9 -1619
rect 161 -1684 178 -1619
rect 230 -1684 247 -1619
rect 301 -1684 318 -1619
rect 446 -1684 463 -1619
rect 616 -1684 633 -1619
rect 685 -1684 702 -1619
rect 756 -1684 773 -1619
rect 901 -1684 918 -1619
rect 1071 -1684 1088 -1619
rect 1140 -1684 1157 -1619
rect 1211 -1684 1228 -1619
rect 1356 -1684 1373 -1619
<< pmos >>
rect -574 -867 -557 -803
rect -437 -867 -420 -803
rect -289 -867 -272 -803
rect -220 -867 -203 -803
rect -149 -867 -132 -803
rect -4 -867 13 -803
rect 163 -867 180 -803
rect 232 -867 249 -803
rect 303 -867 320 -803
rect 448 -867 465 -803
rect 618 -867 635 -803
rect 687 -867 704 -803
rect 758 -867 775 -803
rect 903 -867 920 -803
rect 1068 -867 1085 -803
rect 1137 -867 1154 -803
rect 1208 -867 1225 -803
rect 1353 -867 1370 -803
rect -445 -1419 -428 -1355
rect -293 -1419 -276 -1355
rect -224 -1419 -207 -1355
rect -153 -1419 -136 -1355
rect -8 -1419 9 -1355
rect 161 -1419 178 -1355
rect 230 -1419 247 -1355
rect 301 -1419 318 -1355
rect 446 -1419 463 -1355
rect 616 -1419 633 -1355
rect 685 -1419 702 -1355
rect 756 -1419 773 -1355
rect 901 -1419 918 -1355
rect 1071 -1419 1088 -1355
rect 1140 -1419 1157 -1355
rect 1211 -1419 1228 -1355
rect 1356 -1419 1373 -1355
<< ndiff >>
rect -619 -1079 -574 -1067
rect -619 -1120 -610 -1079
rect -588 -1120 -574 -1079
rect -619 -1132 -574 -1120
rect -557 -1079 -511 -1067
rect -557 -1120 -543 -1079
rect -521 -1120 -511 -1079
rect -557 -1132 -511 -1120
rect -482 -1079 -437 -1067
rect -482 -1120 -473 -1079
rect -451 -1120 -437 -1079
rect -482 -1132 -437 -1120
rect -420 -1079 -374 -1067
rect -420 -1120 -406 -1079
rect -384 -1120 -374 -1079
rect -420 -1132 -374 -1120
rect -336 -1080 -289 -1067
rect -336 -1121 -321 -1080
rect -299 -1121 -289 -1080
rect -336 -1132 -289 -1121
rect -272 -1132 -220 -1067
rect -203 -1132 -149 -1067
rect -132 -1078 -85 -1067
rect -132 -1119 -120 -1078
rect -98 -1119 -85 -1078
rect -132 -1132 -85 -1119
rect -50 -1079 -4 -1067
rect -50 -1120 -40 -1079
rect -18 -1120 -4 -1079
rect -50 -1132 -4 -1120
rect 13 -1079 59 -1067
rect 13 -1120 27 -1079
rect 49 -1120 59 -1079
rect 13 -1132 59 -1120
rect 116 -1080 163 -1067
rect 116 -1121 131 -1080
rect 153 -1121 163 -1080
rect 116 -1132 163 -1121
rect 180 -1132 232 -1067
rect 249 -1132 303 -1067
rect 320 -1078 367 -1067
rect 320 -1119 332 -1078
rect 354 -1119 367 -1078
rect 320 -1132 367 -1119
rect 402 -1079 448 -1067
rect 402 -1120 412 -1079
rect 434 -1120 448 -1079
rect 402 -1132 448 -1120
rect 465 -1079 511 -1067
rect 465 -1120 479 -1079
rect 501 -1120 511 -1079
rect 465 -1132 511 -1120
rect 571 -1080 618 -1067
rect 571 -1121 586 -1080
rect 608 -1121 618 -1080
rect 571 -1132 618 -1121
rect 635 -1132 687 -1067
rect 704 -1132 758 -1067
rect 775 -1078 822 -1067
rect 775 -1119 787 -1078
rect 809 -1119 822 -1078
rect 775 -1132 822 -1119
rect 857 -1079 903 -1067
rect 857 -1120 867 -1079
rect 889 -1120 903 -1079
rect 857 -1132 903 -1120
rect 920 -1079 966 -1067
rect 920 -1120 934 -1079
rect 956 -1120 966 -1079
rect 920 -1132 966 -1120
rect 1021 -1080 1068 -1067
rect 1021 -1121 1036 -1080
rect 1058 -1121 1068 -1080
rect 1021 -1132 1068 -1121
rect 1085 -1132 1137 -1067
rect 1154 -1132 1208 -1067
rect 1225 -1078 1272 -1067
rect 1225 -1119 1237 -1078
rect 1259 -1119 1272 -1078
rect 1225 -1132 1272 -1119
rect 1307 -1079 1353 -1067
rect 1307 -1120 1317 -1079
rect 1339 -1120 1353 -1079
rect 1307 -1132 1353 -1120
rect 1370 -1079 1416 -1067
rect 1370 -1120 1384 -1079
rect 1406 -1120 1416 -1079
rect 1370 -1132 1416 -1120
rect -490 -1631 -445 -1619
rect -490 -1672 -481 -1631
rect -459 -1672 -445 -1631
rect -490 -1684 -445 -1672
rect -428 -1631 -382 -1619
rect -428 -1672 -414 -1631
rect -392 -1672 -382 -1631
rect -428 -1684 -382 -1672
rect -340 -1632 -293 -1619
rect -340 -1673 -325 -1632
rect -303 -1673 -293 -1632
rect -340 -1684 -293 -1673
rect -276 -1684 -224 -1619
rect -207 -1684 -153 -1619
rect -136 -1630 -89 -1619
rect -136 -1671 -124 -1630
rect -102 -1671 -89 -1630
rect -136 -1684 -89 -1671
rect -54 -1631 -8 -1619
rect -54 -1672 -44 -1631
rect -22 -1672 -8 -1631
rect -54 -1684 -8 -1672
rect 9 -1631 55 -1619
rect 9 -1672 23 -1631
rect 45 -1672 55 -1631
rect 9 -1684 55 -1672
rect 114 -1632 161 -1619
rect 114 -1673 129 -1632
rect 151 -1673 161 -1632
rect 114 -1684 161 -1673
rect 178 -1684 230 -1619
rect 247 -1684 301 -1619
rect 318 -1630 365 -1619
rect 318 -1671 330 -1630
rect 352 -1671 365 -1630
rect 318 -1684 365 -1671
rect 400 -1631 446 -1619
rect 400 -1672 410 -1631
rect 432 -1672 446 -1631
rect 400 -1684 446 -1672
rect 463 -1631 509 -1619
rect 463 -1672 477 -1631
rect 499 -1672 509 -1631
rect 463 -1684 509 -1672
rect 569 -1632 616 -1619
rect 569 -1673 584 -1632
rect 606 -1673 616 -1632
rect 569 -1684 616 -1673
rect 633 -1684 685 -1619
rect 702 -1684 756 -1619
rect 773 -1630 820 -1619
rect 773 -1671 785 -1630
rect 807 -1671 820 -1630
rect 773 -1684 820 -1671
rect 855 -1631 901 -1619
rect 855 -1672 865 -1631
rect 887 -1672 901 -1631
rect 855 -1684 901 -1672
rect 918 -1631 964 -1619
rect 918 -1672 932 -1631
rect 954 -1672 964 -1631
rect 918 -1684 964 -1672
rect 1024 -1632 1071 -1619
rect 1024 -1673 1039 -1632
rect 1061 -1673 1071 -1632
rect 1024 -1684 1071 -1673
rect 1088 -1684 1140 -1619
rect 1157 -1684 1211 -1619
rect 1228 -1630 1275 -1619
rect 1228 -1671 1240 -1630
rect 1262 -1671 1275 -1630
rect 1228 -1684 1275 -1671
rect 1310 -1631 1356 -1619
rect 1310 -1672 1320 -1631
rect 1342 -1672 1356 -1631
rect 1310 -1684 1356 -1672
rect 1373 -1631 1419 -1619
rect 1373 -1672 1387 -1631
rect 1409 -1672 1419 -1631
rect 1373 -1684 1419 -1672
<< pdiff >>
rect -619 -819 -574 -803
rect -619 -854 -606 -819
rect -581 -854 -574 -819
rect -619 -867 -574 -854
rect -557 -819 -511 -803
rect -557 -854 -544 -819
rect -519 -854 -511 -819
rect -557 -867 -511 -854
rect -482 -819 -437 -803
rect -482 -854 -469 -819
rect -444 -854 -437 -819
rect -482 -867 -437 -854
rect -420 -819 -374 -803
rect -420 -854 -407 -819
rect -382 -854 -374 -819
rect -420 -867 -374 -854
rect -337 -818 -289 -803
rect -337 -853 -324 -818
rect -299 -853 -289 -818
rect -337 -867 -289 -853
rect -272 -816 -220 -803
rect -272 -851 -258 -816
rect -233 -851 -220 -816
rect -272 -867 -220 -851
rect -203 -817 -149 -803
rect -203 -852 -189 -817
rect -164 -852 -149 -817
rect -203 -867 -149 -852
rect -132 -818 -84 -803
rect -132 -853 -121 -818
rect -96 -853 -84 -818
rect -132 -867 -84 -853
rect -49 -819 -4 -803
rect -49 -854 -36 -819
rect -11 -854 -4 -819
rect -49 -867 -4 -854
rect 13 -819 59 -803
rect 13 -854 26 -819
rect 51 -854 59 -819
rect 13 -867 59 -854
rect 115 -818 163 -803
rect 115 -853 128 -818
rect 153 -853 163 -818
rect 115 -867 163 -853
rect 180 -816 232 -803
rect 180 -851 194 -816
rect 219 -851 232 -816
rect 180 -867 232 -851
rect 249 -817 303 -803
rect 249 -852 263 -817
rect 288 -852 303 -817
rect 249 -867 303 -852
rect 320 -818 368 -803
rect 320 -853 331 -818
rect 356 -853 368 -818
rect 320 -867 368 -853
rect 403 -819 448 -803
rect 403 -854 416 -819
rect 441 -854 448 -819
rect 403 -867 448 -854
rect 465 -819 511 -803
rect 465 -854 478 -819
rect 503 -854 511 -819
rect 465 -867 511 -854
rect 570 -818 618 -803
rect 570 -853 583 -818
rect 608 -853 618 -818
rect 570 -867 618 -853
rect 635 -816 687 -803
rect 635 -851 649 -816
rect 674 -851 687 -816
rect 635 -867 687 -851
rect 704 -817 758 -803
rect 704 -852 718 -817
rect 743 -852 758 -817
rect 704 -867 758 -852
rect 775 -818 823 -803
rect 775 -853 786 -818
rect 811 -853 823 -818
rect 775 -867 823 -853
rect 858 -819 903 -803
rect 858 -854 871 -819
rect 896 -854 903 -819
rect 858 -867 903 -854
rect 920 -819 966 -803
rect 920 -854 933 -819
rect 958 -854 966 -819
rect 920 -867 966 -854
rect 1020 -818 1068 -803
rect 1020 -853 1033 -818
rect 1058 -853 1068 -818
rect 1020 -867 1068 -853
rect 1085 -816 1137 -803
rect 1085 -851 1099 -816
rect 1124 -851 1137 -816
rect 1085 -867 1137 -851
rect 1154 -817 1208 -803
rect 1154 -852 1168 -817
rect 1193 -852 1208 -817
rect 1154 -867 1208 -852
rect 1225 -818 1273 -803
rect 1225 -853 1236 -818
rect 1261 -853 1273 -818
rect 1225 -867 1273 -853
rect 1308 -819 1353 -803
rect 1308 -854 1321 -819
rect 1346 -854 1353 -819
rect 1308 -867 1353 -854
rect 1370 -819 1416 -803
rect 1370 -854 1383 -819
rect 1408 -854 1416 -819
rect 1370 -867 1416 -854
rect -490 -1371 -445 -1355
rect -490 -1406 -477 -1371
rect -452 -1406 -445 -1371
rect -490 -1419 -445 -1406
rect -428 -1371 -382 -1355
rect -428 -1406 -415 -1371
rect -390 -1406 -382 -1371
rect -428 -1419 -382 -1406
rect -341 -1370 -293 -1355
rect -341 -1405 -328 -1370
rect -303 -1405 -293 -1370
rect -341 -1419 -293 -1405
rect -276 -1368 -224 -1355
rect -276 -1403 -262 -1368
rect -237 -1403 -224 -1368
rect -276 -1419 -224 -1403
rect -207 -1369 -153 -1355
rect -207 -1404 -193 -1369
rect -168 -1404 -153 -1369
rect -207 -1419 -153 -1404
rect -136 -1370 -88 -1355
rect -136 -1405 -125 -1370
rect -100 -1405 -88 -1370
rect -136 -1419 -88 -1405
rect -53 -1371 -8 -1355
rect -53 -1406 -40 -1371
rect -15 -1406 -8 -1371
rect -53 -1419 -8 -1406
rect 9 -1371 55 -1355
rect 9 -1406 22 -1371
rect 47 -1406 55 -1371
rect 9 -1419 55 -1406
rect 113 -1370 161 -1355
rect 113 -1405 126 -1370
rect 151 -1405 161 -1370
rect 113 -1419 161 -1405
rect 178 -1368 230 -1355
rect 178 -1403 192 -1368
rect 217 -1403 230 -1368
rect 178 -1419 230 -1403
rect 247 -1369 301 -1355
rect 247 -1404 261 -1369
rect 286 -1404 301 -1369
rect 247 -1419 301 -1404
rect 318 -1370 366 -1355
rect 318 -1405 329 -1370
rect 354 -1405 366 -1370
rect 318 -1419 366 -1405
rect 401 -1371 446 -1355
rect 401 -1406 414 -1371
rect 439 -1406 446 -1371
rect 401 -1419 446 -1406
rect 463 -1371 509 -1355
rect 463 -1406 476 -1371
rect 501 -1406 509 -1371
rect 463 -1419 509 -1406
rect 568 -1370 616 -1355
rect 568 -1405 581 -1370
rect 606 -1405 616 -1370
rect 568 -1419 616 -1405
rect 633 -1368 685 -1355
rect 633 -1403 647 -1368
rect 672 -1403 685 -1368
rect 633 -1419 685 -1403
rect 702 -1369 756 -1355
rect 702 -1404 716 -1369
rect 741 -1404 756 -1369
rect 702 -1419 756 -1404
rect 773 -1370 821 -1355
rect 773 -1405 784 -1370
rect 809 -1405 821 -1370
rect 773 -1419 821 -1405
rect 856 -1371 901 -1355
rect 856 -1406 869 -1371
rect 894 -1406 901 -1371
rect 856 -1419 901 -1406
rect 918 -1371 964 -1355
rect 918 -1406 931 -1371
rect 956 -1406 964 -1371
rect 918 -1419 964 -1406
rect 1023 -1370 1071 -1355
rect 1023 -1405 1036 -1370
rect 1061 -1405 1071 -1370
rect 1023 -1419 1071 -1405
rect 1088 -1368 1140 -1355
rect 1088 -1403 1102 -1368
rect 1127 -1403 1140 -1368
rect 1088 -1419 1140 -1403
rect 1157 -1369 1211 -1355
rect 1157 -1404 1171 -1369
rect 1196 -1404 1211 -1369
rect 1157 -1419 1211 -1404
rect 1228 -1370 1276 -1355
rect 1228 -1405 1239 -1370
rect 1264 -1405 1276 -1370
rect 1228 -1419 1276 -1405
rect 1311 -1371 1356 -1355
rect 1311 -1406 1324 -1371
rect 1349 -1406 1356 -1371
rect 1311 -1419 1356 -1406
rect 1373 -1371 1419 -1355
rect 1373 -1406 1386 -1371
rect 1411 -1406 1419 -1371
rect 1373 -1419 1419 -1406
<< ndiffc >>
rect -610 -1120 -588 -1079
rect -543 -1120 -521 -1079
rect -473 -1120 -451 -1079
rect -406 -1120 -384 -1079
rect -321 -1121 -299 -1080
rect -120 -1119 -98 -1078
rect -40 -1120 -18 -1079
rect 27 -1120 49 -1079
rect 131 -1121 153 -1080
rect 332 -1119 354 -1078
rect 412 -1120 434 -1079
rect 479 -1120 501 -1079
rect 586 -1121 608 -1080
rect 787 -1119 809 -1078
rect 867 -1120 889 -1079
rect 934 -1120 956 -1079
rect 1036 -1121 1058 -1080
rect 1237 -1119 1259 -1078
rect 1317 -1120 1339 -1079
rect 1384 -1120 1406 -1079
rect -481 -1672 -459 -1631
rect -414 -1672 -392 -1631
rect -325 -1673 -303 -1632
rect -124 -1671 -102 -1630
rect -44 -1672 -22 -1631
rect 23 -1672 45 -1631
rect 129 -1673 151 -1632
rect 330 -1671 352 -1630
rect 410 -1672 432 -1631
rect 477 -1672 499 -1631
rect 584 -1673 606 -1632
rect 785 -1671 807 -1630
rect 865 -1672 887 -1631
rect 932 -1672 954 -1631
rect 1039 -1673 1061 -1632
rect 1240 -1671 1262 -1630
rect 1320 -1672 1342 -1631
rect 1387 -1672 1409 -1631
<< pdiffc >>
rect -606 -854 -581 -819
rect -544 -854 -519 -819
rect -469 -854 -444 -819
rect -407 -854 -382 -819
rect -324 -853 -299 -818
rect -258 -851 -233 -816
rect -189 -852 -164 -817
rect -121 -853 -96 -818
rect -36 -854 -11 -819
rect 26 -854 51 -819
rect 128 -853 153 -818
rect 194 -851 219 -816
rect 263 -852 288 -817
rect 331 -853 356 -818
rect 416 -854 441 -819
rect 478 -854 503 -819
rect 583 -853 608 -818
rect 649 -851 674 -816
rect 718 -852 743 -817
rect 786 -853 811 -818
rect 871 -854 896 -819
rect 933 -854 958 -819
rect 1033 -853 1058 -818
rect 1099 -851 1124 -816
rect 1168 -852 1193 -817
rect 1236 -853 1261 -818
rect 1321 -854 1346 -819
rect 1383 -854 1408 -819
rect -477 -1406 -452 -1371
rect -415 -1406 -390 -1371
rect -328 -1405 -303 -1370
rect -262 -1403 -237 -1368
rect -193 -1404 -168 -1369
rect -125 -1405 -100 -1370
rect -40 -1406 -15 -1371
rect 22 -1406 47 -1371
rect 126 -1405 151 -1370
rect 192 -1403 217 -1368
rect 261 -1404 286 -1369
rect 329 -1405 354 -1370
rect 414 -1406 439 -1371
rect 476 -1406 501 -1371
rect 581 -1405 606 -1370
rect 647 -1403 672 -1368
rect 716 -1404 741 -1369
rect 784 -1405 809 -1370
rect 869 -1406 894 -1371
rect 931 -1406 956 -1371
rect 1036 -1405 1061 -1370
rect 1102 -1403 1127 -1368
rect 1171 -1404 1196 -1369
rect 1239 -1405 1264 -1370
rect 1324 -1406 1349 -1371
rect 1386 -1406 1411 -1371
<< psubdiff >>
rect -619 -1186 1437 -1181
rect -619 -1187 -290 -1186
rect -619 -1208 -575 -1187
rect -554 -1208 -534 -1187
rect -513 -1208 -438 -1187
rect -417 -1208 -397 -1187
rect -376 -1207 -290 -1187
rect -269 -1187 -203 -1186
rect -269 -1207 -247 -1187
rect -376 -1208 -247 -1207
rect -226 -1207 -203 -1187
rect -182 -1207 -159 -1186
rect -138 -1187 162 -1186
rect -138 -1207 -119 -1187
rect -226 -1208 -119 -1207
rect -98 -1208 -75 -1187
rect -54 -1208 -5 -1187
rect 16 -1208 36 -1187
rect 57 -1207 162 -1187
rect 183 -1187 249 -1186
rect 183 -1207 205 -1187
rect 57 -1208 205 -1207
rect 226 -1207 249 -1187
rect 270 -1207 293 -1186
rect 314 -1187 617 -1186
rect 314 -1207 333 -1187
rect 226 -1208 333 -1207
rect 354 -1208 377 -1187
rect 398 -1208 447 -1187
rect 468 -1208 488 -1187
rect 509 -1207 617 -1187
rect 638 -1187 704 -1186
rect 638 -1207 660 -1187
rect 509 -1208 660 -1207
rect 681 -1207 704 -1187
rect 725 -1207 748 -1186
rect 769 -1187 1067 -1186
rect 769 -1207 788 -1187
rect 681 -1208 788 -1207
rect 809 -1208 832 -1187
rect 853 -1208 902 -1187
rect 923 -1208 943 -1187
rect 964 -1207 1067 -1187
rect 1088 -1187 1154 -1186
rect 1088 -1207 1110 -1187
rect 964 -1208 1110 -1207
rect 1131 -1207 1154 -1187
rect 1175 -1207 1198 -1186
rect 1219 -1187 1437 -1186
rect 1219 -1207 1238 -1187
rect 1131 -1208 1238 -1207
rect 1259 -1208 1282 -1187
rect 1303 -1208 1352 -1187
rect 1373 -1208 1393 -1187
rect 1414 -1208 1437 -1187
rect -619 -1216 1437 -1208
rect -490 -1738 1452 -1733
rect -490 -1739 -294 -1738
rect -490 -1760 -446 -1739
rect -425 -1760 -405 -1739
rect -384 -1759 -294 -1739
rect -273 -1739 -207 -1738
rect -273 -1759 -251 -1739
rect -384 -1760 -251 -1759
rect -230 -1759 -207 -1739
rect -186 -1759 -163 -1738
rect -142 -1739 160 -1738
rect -142 -1759 -123 -1739
rect -230 -1760 -123 -1759
rect -102 -1760 -79 -1739
rect -58 -1760 -9 -1739
rect 12 -1760 32 -1739
rect 53 -1759 160 -1739
rect 181 -1739 247 -1738
rect 181 -1759 203 -1739
rect 53 -1760 203 -1759
rect 224 -1759 247 -1739
rect 268 -1759 291 -1738
rect 312 -1739 615 -1738
rect 312 -1759 331 -1739
rect 224 -1760 331 -1759
rect 352 -1760 375 -1739
rect 396 -1760 445 -1739
rect 466 -1760 486 -1739
rect 507 -1759 615 -1739
rect 636 -1739 702 -1738
rect 636 -1759 658 -1739
rect 507 -1760 658 -1759
rect 679 -1759 702 -1739
rect 723 -1759 746 -1738
rect 767 -1739 1070 -1738
rect 767 -1759 786 -1739
rect 679 -1760 786 -1759
rect 807 -1760 830 -1739
rect 851 -1760 900 -1739
rect 921 -1760 941 -1739
rect 962 -1759 1070 -1739
rect 1091 -1739 1157 -1738
rect 1091 -1759 1113 -1739
rect 962 -1760 1113 -1759
rect 1134 -1759 1157 -1739
rect 1178 -1759 1201 -1738
rect 1222 -1739 1452 -1738
rect 1222 -1759 1241 -1739
rect 1134 -1760 1241 -1759
rect 1262 -1760 1285 -1739
rect 1306 -1760 1355 -1739
rect 1376 -1760 1396 -1739
rect 1417 -1760 1452 -1739
rect -490 -1768 1452 -1760
<< nsubdiff >>
rect -619 -703 79 -699
rect -619 -705 -84 -703
rect -619 -726 -563 -705
rect -542 -706 -426 -705
rect -542 -726 -524 -706
rect -619 -727 -524 -726
rect -503 -726 -426 -706
rect -405 -706 -276 -705
rect -405 -726 -387 -706
rect -503 -727 -387 -726
rect -366 -726 -276 -706
rect -255 -706 -141 -705
rect -255 -726 -232 -706
rect -366 -727 -232 -726
rect -211 -726 -141 -706
rect -120 -724 -84 -705
rect -63 -705 79 -703
rect -63 -724 7 -705
rect -120 -726 7 -724
rect 28 -706 79 -705
rect 28 -726 46 -706
rect -211 -727 46 -726
rect 67 -727 79 -706
rect -619 -734 79 -727
rect 114 -703 531 -699
rect 114 -705 368 -703
rect 114 -726 176 -705
rect 197 -706 311 -705
rect 197 -726 220 -706
rect 114 -727 220 -726
rect 241 -726 311 -706
rect 332 -724 368 -705
rect 389 -705 531 -703
rect 389 -724 459 -705
rect 332 -726 459 -724
rect 480 -706 531 -705
rect 480 -726 498 -706
rect 241 -727 498 -726
rect 519 -727 531 -706
rect 114 -734 531 -727
rect 569 -703 986 -699
rect 569 -705 823 -703
rect 569 -726 631 -705
rect 652 -706 766 -705
rect 652 -726 675 -706
rect 569 -727 675 -726
rect 696 -726 766 -706
rect 787 -724 823 -705
rect 844 -705 986 -703
rect 844 -724 914 -705
rect 787 -726 914 -724
rect 935 -706 986 -705
rect 935 -726 953 -706
rect 696 -727 953 -726
rect 974 -727 986 -706
rect 569 -734 986 -727
rect 1019 -703 1419 -699
rect 1019 -705 1273 -703
rect 1019 -726 1081 -705
rect 1102 -706 1216 -705
rect 1102 -726 1125 -706
rect 1019 -727 1125 -726
rect 1146 -726 1216 -706
rect 1237 -724 1273 -705
rect 1294 -705 1419 -703
rect 1294 -724 1364 -705
rect 1237 -726 1364 -724
rect 1385 -726 1419 -705
rect 1146 -727 1419 -726
rect 1019 -734 1419 -727
rect -360 -735 -280 -734
rect -490 -1255 75 -1251
rect -490 -1257 -88 -1255
rect -490 -1278 -434 -1257
rect -413 -1258 -280 -1257
rect -413 -1278 -395 -1258
rect -490 -1279 -395 -1278
rect -374 -1278 -280 -1258
rect -259 -1258 -145 -1257
rect -259 -1278 -236 -1258
rect -374 -1279 -236 -1278
rect -215 -1278 -145 -1258
rect -124 -1276 -88 -1257
rect -67 -1257 75 -1255
rect -67 -1276 3 -1257
rect -124 -1278 3 -1276
rect 24 -1258 75 -1257
rect 24 -1278 42 -1258
rect -215 -1279 42 -1278
rect 63 -1279 75 -1258
rect -490 -1286 75 -1279
rect 112 -1255 529 -1251
rect 112 -1257 366 -1255
rect 112 -1278 174 -1257
rect 195 -1258 309 -1257
rect 195 -1278 218 -1258
rect 112 -1279 218 -1278
rect 239 -1278 309 -1258
rect 330 -1276 366 -1257
rect 387 -1257 529 -1255
rect 387 -1276 457 -1257
rect 330 -1278 457 -1276
rect 478 -1258 529 -1257
rect 478 -1278 496 -1258
rect 239 -1279 496 -1278
rect 517 -1279 529 -1258
rect 112 -1286 529 -1279
rect 567 -1255 984 -1251
rect 567 -1257 821 -1255
rect 567 -1278 629 -1257
rect 650 -1258 764 -1257
rect 650 -1278 673 -1258
rect 567 -1279 673 -1278
rect 694 -1278 764 -1258
rect 785 -1276 821 -1257
rect 842 -1257 984 -1255
rect 842 -1276 912 -1257
rect 785 -1278 912 -1276
rect 933 -1258 984 -1257
rect 933 -1278 951 -1258
rect 694 -1279 951 -1278
rect 972 -1279 984 -1258
rect 567 -1286 984 -1279
rect 1022 -1255 1439 -1251
rect 1022 -1257 1276 -1255
rect 1022 -1278 1084 -1257
rect 1105 -1258 1219 -1257
rect 1105 -1278 1128 -1258
rect 1022 -1279 1128 -1278
rect 1149 -1278 1219 -1258
rect 1240 -1276 1276 -1257
rect 1297 -1257 1439 -1255
rect 1297 -1276 1367 -1257
rect 1240 -1278 1367 -1276
rect 1388 -1258 1439 -1257
rect 1388 -1278 1406 -1258
rect 1149 -1279 1406 -1278
rect 1427 -1279 1439 -1258
rect 1022 -1286 1439 -1279
<< psubdiffcont >>
rect -575 -1208 -554 -1187
rect -534 -1208 -513 -1187
rect -438 -1208 -417 -1187
rect -397 -1208 -376 -1187
rect -290 -1207 -269 -1186
rect -247 -1208 -226 -1187
rect -203 -1207 -182 -1186
rect -159 -1207 -138 -1186
rect -119 -1208 -98 -1187
rect -75 -1208 -54 -1187
rect -5 -1208 16 -1187
rect 36 -1208 57 -1187
rect 162 -1207 183 -1186
rect 205 -1208 226 -1187
rect 249 -1207 270 -1186
rect 293 -1207 314 -1186
rect 333 -1208 354 -1187
rect 377 -1208 398 -1187
rect 447 -1208 468 -1187
rect 488 -1208 509 -1187
rect 617 -1207 638 -1186
rect 660 -1208 681 -1187
rect 704 -1207 725 -1186
rect 748 -1207 769 -1186
rect 788 -1208 809 -1187
rect 832 -1208 853 -1187
rect 902 -1208 923 -1187
rect 943 -1208 964 -1187
rect 1067 -1207 1088 -1186
rect 1110 -1208 1131 -1187
rect 1154 -1207 1175 -1186
rect 1198 -1207 1219 -1186
rect 1238 -1208 1259 -1187
rect 1282 -1208 1303 -1187
rect 1352 -1208 1373 -1187
rect 1393 -1208 1414 -1187
rect -446 -1760 -425 -1739
rect -405 -1760 -384 -1739
rect -294 -1759 -273 -1738
rect -251 -1760 -230 -1739
rect -207 -1759 -186 -1738
rect -163 -1759 -142 -1738
rect -123 -1760 -102 -1739
rect -79 -1760 -58 -1739
rect -9 -1760 12 -1739
rect 32 -1760 53 -1739
rect 160 -1759 181 -1738
rect 203 -1760 224 -1739
rect 247 -1759 268 -1738
rect 291 -1759 312 -1738
rect 331 -1760 352 -1739
rect 375 -1760 396 -1739
rect 445 -1760 466 -1739
rect 486 -1760 507 -1739
rect 615 -1759 636 -1738
rect 658 -1760 679 -1739
rect 702 -1759 723 -1738
rect 746 -1759 767 -1738
rect 786 -1760 807 -1739
rect 830 -1760 851 -1739
rect 900 -1760 921 -1739
rect 941 -1760 962 -1739
rect 1070 -1759 1091 -1738
rect 1113 -1760 1134 -1739
rect 1157 -1759 1178 -1738
rect 1201 -1759 1222 -1738
rect 1241 -1760 1262 -1739
rect 1285 -1760 1306 -1739
rect 1355 -1760 1376 -1739
rect 1396 -1760 1417 -1739
<< nsubdiffcont >>
rect -563 -726 -542 -705
rect -524 -727 -503 -706
rect -426 -726 -405 -705
rect -387 -727 -366 -706
rect -276 -726 -255 -705
rect -232 -727 -211 -706
rect -141 -726 -120 -705
rect -84 -724 -63 -703
rect 7 -726 28 -705
rect 46 -727 67 -706
rect 176 -726 197 -705
rect 220 -727 241 -706
rect 311 -726 332 -705
rect 368 -724 389 -703
rect 459 -726 480 -705
rect 498 -727 519 -706
rect 631 -726 652 -705
rect 675 -727 696 -706
rect 766 -726 787 -705
rect 823 -724 844 -703
rect 914 -726 935 -705
rect 953 -727 974 -706
rect 1081 -726 1102 -705
rect 1125 -727 1146 -706
rect 1216 -726 1237 -705
rect 1273 -724 1294 -703
rect 1364 -726 1385 -705
rect -434 -1278 -413 -1257
rect -395 -1279 -374 -1258
rect -280 -1278 -259 -1257
rect -236 -1279 -215 -1258
rect -145 -1278 -124 -1257
rect -88 -1276 -67 -1255
rect 3 -1278 24 -1257
rect 42 -1279 63 -1258
rect 174 -1278 195 -1257
rect 218 -1279 239 -1258
rect 309 -1278 330 -1257
rect 366 -1276 387 -1255
rect 457 -1278 478 -1257
rect 496 -1279 517 -1258
rect 629 -1278 650 -1257
rect 673 -1279 694 -1258
rect 764 -1278 785 -1257
rect 821 -1276 842 -1255
rect 912 -1278 933 -1257
rect 951 -1279 972 -1258
rect 1084 -1278 1105 -1257
rect 1128 -1279 1149 -1258
rect 1219 -1278 1240 -1257
rect 1276 -1276 1297 -1255
rect 1367 -1278 1388 -1257
rect 1406 -1279 1427 -1258
<< poly >>
rect -574 -803 -557 -771
rect -437 -803 -420 -771
rect -289 -803 -272 -770
rect -220 -803 -203 -770
rect -149 -803 -132 -771
rect -4 -803 13 -771
rect 163 -803 180 -770
rect 232 -803 249 -770
rect 303 -803 320 -771
rect 448 -803 465 -771
rect 618 -803 635 -770
rect 687 -803 704 -770
rect 758 -803 775 -771
rect 903 -803 920 -771
rect 1068 -803 1085 -770
rect 1137 -803 1154 -770
rect 1208 -803 1225 -771
rect 1353 -803 1370 -771
rect -648 -963 -610 -957
rect -574 -963 -557 -867
rect -648 -965 -557 -963
rect -648 -982 -638 -965
rect -621 -978 -557 -965
rect -621 -982 -610 -978
rect -648 -990 -610 -982
rect -574 -1067 -557 -978
rect -437 -980 -420 -867
rect -289 -884 -272 -867
rect -314 -892 -272 -884
rect -314 -913 -304 -892
rect -283 -913 -272 -892
rect -314 -922 -272 -913
rect -468 -989 -420 -980
rect -468 -1011 -456 -989
rect -431 -1011 -420 -989
rect -468 -1022 -420 -1011
rect -437 -1067 -420 -1022
rect -289 -1067 -272 -922
rect -220 -940 -203 -867
rect -242 -949 -201 -940
rect -242 -970 -230 -949
rect -209 -970 -201 -949
rect -242 -978 -201 -970
rect -220 -1067 -203 -978
rect -149 -1002 -132 -867
rect -4 -991 13 -867
rect 163 -884 180 -867
rect 138 -892 180 -884
rect 138 -913 148 -892
rect 169 -913 180 -892
rect 138 -922 180 -913
rect -171 -1009 -132 -1002
rect -171 -1030 -161 -1009
rect -140 -1030 -132 -1009
rect -36 -1000 13 -991
rect -36 -1021 -27 -1000
rect -4 -1021 13 -1000
rect -36 -1029 13 -1021
rect -171 -1040 -132 -1030
rect -149 -1067 -132 -1040
rect -4 -1067 13 -1029
rect 163 -1067 180 -922
rect 232 -940 249 -867
rect 210 -949 251 -940
rect 210 -970 222 -949
rect 243 -970 251 -949
rect 210 -978 251 -970
rect 232 -1067 249 -978
rect 303 -1002 320 -867
rect 350 -949 388 -942
rect 448 -949 465 -867
rect 618 -884 635 -867
rect 593 -892 635 -884
rect 593 -913 603 -892
rect 624 -913 635 -892
rect 593 -922 635 -913
rect 350 -950 465 -949
rect 350 -967 359 -950
rect 377 -964 465 -950
rect 377 -967 388 -964
rect 350 -977 388 -967
rect 281 -1009 320 -1002
rect 281 -1030 291 -1009
rect 312 -1030 320 -1009
rect 281 -1040 320 -1030
rect 303 -1067 320 -1040
rect 448 -1067 465 -964
rect 618 -1067 635 -922
rect 687 -940 704 -867
rect 665 -949 706 -940
rect 665 -970 677 -949
rect 698 -970 706 -949
rect 665 -978 706 -970
rect 687 -1067 704 -978
rect 758 -1002 775 -867
rect 903 -910 920 -867
rect 1068 -884 1085 -867
rect 877 -920 920 -910
rect 877 -938 889 -920
rect 907 -938 920 -920
rect 1043 -892 1085 -884
rect 1043 -913 1053 -892
rect 1074 -913 1085 -892
rect 1043 -922 1085 -913
rect 877 -946 920 -938
rect 736 -1009 775 -1002
rect 736 -1030 746 -1009
rect 767 -1030 775 -1009
rect 736 -1040 775 -1030
rect 758 -1067 775 -1040
rect 903 -1067 920 -946
rect 1068 -1067 1085 -922
rect 1137 -940 1154 -867
rect 1115 -949 1156 -940
rect 1115 -970 1127 -949
rect 1148 -970 1156 -949
rect 1115 -978 1156 -970
rect 1137 -1067 1154 -978
rect 1208 -1002 1225 -867
rect 1353 -950 1370 -867
rect 1320 -958 1370 -950
rect 1320 -976 1330 -958
rect 1348 -976 1370 -958
rect 1320 -986 1370 -976
rect 1186 -1009 1225 -1002
rect 1186 -1030 1196 -1009
rect 1217 -1030 1225 -1009
rect 1186 -1040 1225 -1030
rect 1208 -1067 1225 -1040
rect 1353 -1067 1370 -986
rect -574 -1160 -557 -1132
rect -437 -1160 -420 -1132
rect -289 -1159 -272 -1132
rect -220 -1159 -203 -1132
rect -149 -1160 -132 -1132
rect -4 -1160 13 -1132
rect 163 -1159 180 -1132
rect 232 -1159 249 -1132
rect 303 -1160 320 -1132
rect 448 -1160 465 -1132
rect 618 -1159 635 -1132
rect 687 -1159 704 -1132
rect 758 -1160 775 -1132
rect 903 -1160 920 -1132
rect 1068 -1159 1085 -1132
rect 1137 -1159 1154 -1132
rect 1208 -1160 1225 -1132
rect 1353 -1160 1370 -1132
rect -247 -1309 -206 -1303
rect -445 -1355 -428 -1323
rect -293 -1355 -276 -1322
rect -247 -1329 -239 -1309
rect -217 -1329 -206 -1309
rect -247 -1344 -206 -1329
rect -224 -1355 -207 -1344
rect -153 -1355 -136 -1323
rect -8 -1355 9 -1323
rect 161 -1355 178 -1322
rect 230 -1355 247 -1322
rect 301 -1355 318 -1323
rect 446 -1355 463 -1323
rect 616 -1355 633 -1322
rect 685 -1355 702 -1322
rect 756 -1355 773 -1323
rect 901 -1355 918 -1323
rect 1071 -1355 1088 -1322
rect 1140 -1355 1157 -1322
rect 1211 -1355 1228 -1323
rect 1356 -1355 1373 -1323
rect -445 -1555 -428 -1419
rect -293 -1436 -276 -1419
rect -318 -1444 -276 -1436
rect -318 -1465 -308 -1444
rect -287 -1465 -276 -1444
rect -318 -1474 -276 -1465
rect -463 -1564 -428 -1555
rect -463 -1581 -454 -1564
rect -437 -1581 -428 -1564
rect -463 -1589 -428 -1581
rect -445 -1619 -428 -1589
rect -293 -1619 -276 -1474
rect -224 -1619 -207 -1419
rect -153 -1554 -136 -1419
rect -175 -1561 -136 -1554
rect -175 -1582 -165 -1561
rect -144 -1582 -136 -1561
rect -8 -1569 9 -1419
rect 161 -1436 178 -1419
rect 136 -1444 178 -1436
rect 136 -1465 146 -1444
rect 167 -1465 178 -1444
rect 136 -1474 178 -1465
rect -175 -1592 -136 -1582
rect -153 -1619 -136 -1592
rect -31 -1574 9 -1569
rect -31 -1591 -23 -1574
rect -6 -1591 9 -1574
rect -31 -1599 9 -1591
rect -8 -1619 9 -1599
rect 161 -1619 178 -1474
rect 230 -1492 247 -1419
rect 208 -1501 249 -1492
rect 208 -1522 220 -1501
rect 241 -1522 249 -1501
rect 208 -1530 249 -1522
rect 230 -1619 247 -1530
rect 301 -1554 318 -1419
rect 279 -1561 318 -1554
rect 446 -1555 463 -1419
rect 616 -1436 633 -1419
rect 591 -1444 633 -1436
rect 591 -1465 601 -1444
rect 622 -1465 633 -1444
rect 591 -1474 633 -1465
rect 279 -1582 289 -1561
rect 310 -1582 318 -1561
rect 279 -1592 318 -1582
rect 417 -1564 463 -1555
rect 417 -1581 425 -1564
rect 443 -1581 463 -1564
rect 417 -1588 463 -1581
rect 301 -1619 318 -1592
rect 446 -1619 463 -1588
rect 616 -1619 633 -1474
rect 685 -1492 702 -1419
rect 663 -1501 704 -1492
rect 663 -1522 675 -1501
rect 696 -1522 704 -1501
rect 663 -1530 704 -1522
rect 685 -1619 702 -1530
rect 756 -1554 773 -1419
rect 730 -1563 773 -1554
rect 901 -1557 918 -1419
rect 1071 -1436 1088 -1419
rect 1046 -1444 1088 -1436
rect 1046 -1465 1056 -1444
rect 1077 -1465 1088 -1444
rect 1046 -1474 1088 -1465
rect 730 -1584 740 -1563
rect 765 -1584 773 -1563
rect 730 -1593 773 -1584
rect 874 -1564 918 -1557
rect 874 -1582 882 -1564
rect 900 -1582 918 -1564
rect 874 -1590 918 -1582
rect 756 -1619 773 -1593
rect 901 -1619 918 -1590
rect 1071 -1619 1088 -1474
rect 1140 -1492 1157 -1419
rect 1118 -1501 1159 -1492
rect 1118 -1522 1130 -1501
rect 1151 -1522 1159 -1501
rect 1118 -1530 1159 -1522
rect 1140 -1619 1157 -1530
rect 1211 -1554 1228 -1419
rect 1189 -1561 1228 -1554
rect 1356 -1557 1373 -1419
rect 1189 -1582 1199 -1561
rect 1220 -1582 1228 -1561
rect 1189 -1592 1228 -1582
rect 1326 -1565 1373 -1557
rect 1326 -1583 1335 -1565
rect 1353 -1583 1373 -1565
rect 1326 -1591 1373 -1583
rect 1211 -1619 1228 -1592
rect 1356 -1619 1373 -1591
rect -445 -1712 -428 -1684
rect -293 -1711 -276 -1684
rect -224 -1711 -207 -1684
rect -153 -1712 -136 -1684
rect -8 -1712 9 -1684
rect 161 -1711 178 -1684
rect 230 -1711 247 -1684
rect 301 -1712 318 -1684
rect 446 -1712 463 -1684
rect 616 -1711 633 -1684
rect 685 -1711 702 -1684
rect 756 -1712 773 -1684
rect 901 -1712 918 -1684
rect 1071 -1711 1088 -1684
rect 1140 -1711 1157 -1684
rect 1211 -1712 1228 -1684
rect 1356 -1712 1373 -1684
<< polycont >>
rect -638 -982 -621 -965
rect -304 -913 -283 -892
rect -456 -1011 -431 -989
rect -230 -970 -209 -949
rect 148 -913 169 -892
rect -161 -1030 -140 -1009
rect -27 -1021 -4 -1000
rect 222 -970 243 -949
rect 603 -913 624 -892
rect 359 -967 377 -950
rect 291 -1030 312 -1009
rect 677 -970 698 -949
rect 889 -938 907 -920
rect 1053 -913 1074 -892
rect 746 -1030 767 -1009
rect 1127 -970 1148 -949
rect 1330 -976 1348 -958
rect 1196 -1030 1217 -1009
rect -239 -1329 -217 -1309
rect -308 -1465 -287 -1444
rect -454 -1581 -437 -1564
rect -165 -1582 -144 -1561
rect 146 -1465 167 -1444
rect -23 -1591 -6 -1574
rect 220 -1522 241 -1501
rect 601 -1465 622 -1444
rect 289 -1582 310 -1561
rect 425 -1581 443 -1564
rect 675 -1522 696 -1501
rect 1056 -1465 1077 -1444
rect 740 -1584 765 -1563
rect 882 -1582 900 -1564
rect 1130 -1522 1151 -1501
rect 1199 -1582 1220 -1561
rect 1335 -1583 1353 -1565
<< locali >>
rect -619 -703 1437 -699
rect -619 -705 -84 -703
rect -619 -726 -605 -705
rect -584 -726 -563 -705
rect -542 -706 -468 -705
rect -542 -726 -524 -706
rect -619 -727 -524 -726
rect -503 -726 -468 -706
rect -447 -726 -426 -705
rect -405 -706 -319 -705
rect -405 -726 -387 -706
rect -503 -727 -387 -726
rect -366 -726 -319 -706
rect -298 -726 -276 -705
rect -255 -706 -141 -705
rect -255 -726 -232 -706
rect -366 -727 -232 -726
rect -211 -727 -187 -706
rect -166 -726 -141 -706
rect -120 -724 -84 -705
rect -63 -705 368 -703
rect -63 -724 -35 -705
rect -120 -726 -35 -724
rect -14 -726 7 -705
rect 28 -706 133 -705
rect 28 -726 46 -706
rect -166 -727 46 -726
rect 67 -726 133 -706
rect 154 -726 176 -705
rect 197 -706 311 -705
rect 197 -726 220 -706
rect 67 -727 220 -726
rect 241 -727 265 -706
rect 286 -726 311 -706
rect 332 -724 368 -705
rect 389 -705 823 -703
rect 389 -724 417 -705
rect 332 -726 417 -724
rect 438 -726 459 -705
rect 480 -706 588 -705
rect 480 -726 498 -706
rect 286 -727 498 -726
rect 519 -726 588 -706
rect 609 -726 631 -705
rect 652 -706 766 -705
rect 652 -726 675 -706
rect 519 -727 675 -726
rect 696 -727 720 -706
rect 741 -726 766 -706
rect 787 -724 823 -705
rect 844 -705 1273 -703
rect 844 -724 872 -705
rect 787 -726 872 -724
rect 893 -726 914 -705
rect 935 -706 1038 -705
rect 935 -726 953 -706
rect 741 -727 953 -726
rect 974 -726 1038 -706
rect 1059 -726 1081 -705
rect 1102 -706 1216 -705
rect 1102 -726 1125 -706
rect 974 -727 1125 -726
rect 1146 -727 1170 -706
rect 1191 -726 1216 -706
rect 1237 -724 1273 -705
rect 1294 -705 1437 -703
rect 1294 -724 1322 -705
rect 1237 -726 1322 -724
rect 1343 -726 1364 -705
rect 1385 -726 1437 -705
rect 1191 -727 1437 -726
rect -619 -734 1437 -727
rect -605 -803 -584 -734
rect -468 -803 -447 -734
rect -322 -803 -297 -734
rect -188 -803 -163 -734
rect -35 -803 -14 -734
rect 130 -803 155 -734
rect 264 -803 289 -734
rect 417 -803 438 -734
rect 585 -803 610 -734
rect 719 -803 744 -734
rect 872 -803 893 -734
rect 1035 -803 1060 -734
rect 1169 -803 1194 -734
rect 1322 -803 1343 -734
rect -619 -819 -575 -803
rect -619 -854 -606 -819
rect -581 -854 -575 -819
rect -619 -867 -575 -854
rect -556 -819 -511 -803
rect -556 -854 -544 -819
rect -519 -854 -511 -819
rect -556 -867 -511 -854
rect -482 -819 -438 -803
rect -482 -854 -469 -819
rect -444 -854 -438 -819
rect -482 -867 -438 -854
rect -419 -819 -374 -803
rect -419 -854 -407 -819
rect -382 -854 -374 -819
rect -419 -867 -374 -854
rect -337 -818 -290 -803
rect -337 -853 -324 -818
rect -299 -853 -290 -818
rect -337 -867 -290 -853
rect -271 -816 -221 -803
rect -271 -851 -258 -816
rect -233 -851 -221 -816
rect -271 -867 -221 -851
rect -202 -817 -150 -803
rect -202 -852 -189 -817
rect -164 -852 -150 -817
rect -202 -867 -150 -852
rect -131 -818 -84 -803
rect -131 -853 -121 -818
rect -96 -853 -84 -818
rect -131 -867 -84 -853
rect -49 -819 -5 -803
rect -49 -854 -36 -819
rect -11 -854 -5 -819
rect -49 -867 -5 -854
rect 14 -819 59 -803
rect 14 -854 26 -819
rect 51 -854 59 -819
rect 14 -867 59 -854
rect 115 -818 162 -803
rect 115 -853 128 -818
rect 153 -853 162 -818
rect 115 -867 162 -853
rect 181 -816 231 -803
rect 181 -851 194 -816
rect 219 -851 231 -816
rect 181 -867 231 -851
rect 250 -817 302 -803
rect 250 -852 263 -817
rect 288 -852 302 -817
rect 250 -867 302 -852
rect 321 -818 368 -803
rect 321 -853 331 -818
rect 356 -853 368 -818
rect 321 -867 368 -853
rect 403 -819 447 -803
rect 403 -854 416 -819
rect 441 -854 447 -819
rect 403 -867 447 -854
rect 466 -819 511 -803
rect 466 -854 478 -819
rect 503 -854 511 -819
rect 466 -867 511 -854
rect 570 -818 617 -803
rect 570 -853 583 -818
rect 608 -853 617 -818
rect 570 -867 617 -853
rect 636 -816 686 -803
rect 636 -851 649 -816
rect 674 -851 686 -816
rect 636 -867 686 -851
rect 705 -817 757 -803
rect 705 -852 718 -817
rect 743 -852 757 -817
rect 705 -867 757 -852
rect 776 -818 823 -803
rect 776 -853 786 -818
rect 811 -853 823 -818
rect 776 -867 823 -853
rect 858 -819 902 -803
rect 858 -854 871 -819
rect 896 -854 902 -819
rect 858 -867 902 -854
rect 921 -819 966 -803
rect 921 -854 933 -819
rect 958 -854 966 -819
rect 921 -867 966 -854
rect 1020 -818 1067 -803
rect 1020 -853 1033 -818
rect 1058 -853 1067 -818
rect 1020 -867 1067 -853
rect 1086 -816 1136 -803
rect 1086 -851 1099 -816
rect 1124 -851 1136 -816
rect 1086 -867 1136 -851
rect 1155 -817 1207 -803
rect 1155 -852 1168 -817
rect 1193 -852 1207 -817
rect 1155 -867 1207 -852
rect 1226 -818 1273 -803
rect 1226 -853 1236 -818
rect 1261 -853 1273 -818
rect 1226 -867 1273 -853
rect 1308 -819 1352 -803
rect 1308 -854 1321 -819
rect 1346 -854 1352 -819
rect 1308 -867 1352 -854
rect 1371 -819 1416 -803
rect 1371 -854 1383 -819
rect 1408 -854 1416 -819
rect 1371 -867 1416 -854
rect -543 -885 -522 -867
rect -543 -895 -500 -885
rect -543 -912 -530 -895
rect -511 -912 -500 -895
rect -543 -923 -500 -912
rect -648 -965 -610 -957
rect -648 -982 -638 -965
rect -621 -982 -610 -965
rect -648 -990 -610 -982
rect -543 -1067 -522 -923
rect -406 -953 -385 -867
rect -256 -884 -239 -867
rect -102 -884 -85 -867
rect -314 -892 -273 -884
rect -314 -913 -304 -892
rect -283 -913 -273 -892
rect -256 -902 -85 -884
rect -314 -922 -273 -913
rect -242 -949 -201 -940
rect -242 -953 -230 -949
rect -406 -970 -230 -953
rect -209 -970 -201 -949
rect -406 -971 -201 -970
rect -468 -989 -423 -980
rect -468 -1011 -456 -989
rect -431 -1011 -423 -989
rect -468 -1022 -423 -1011
rect -406 -1067 -385 -971
rect -242 -978 -201 -971
rect -171 -1009 -132 -1002
rect -171 -1030 -161 -1009
rect -140 -1030 -132 -1009
rect -171 -1040 -132 -1030
rect -102 -1003 -85 -902
rect -36 -1000 3 -991
rect -36 -1003 -27 -1000
rect -102 -1020 -27 -1003
rect -102 -1067 -85 -1020
rect -36 -1021 -27 -1020
rect -4 -1021 3 -1000
rect -36 -1029 3 -1021
rect 27 -1067 48 -867
rect 196 -884 213 -867
rect 350 -884 367 -867
rect 138 -892 179 -884
rect 138 -913 148 -892
rect 169 -913 179 -892
rect 196 -902 367 -884
rect 138 -922 179 -913
rect 210 -949 251 -940
rect 210 -970 222 -949
rect 243 -970 251 -949
rect 210 -978 251 -970
rect 350 -942 367 -902
rect 350 -950 388 -942
rect 350 -967 359 -950
rect 377 -967 388 -950
rect 350 -977 388 -967
rect 281 -1009 320 -1002
rect 281 -1030 291 -1009
rect 312 -1030 320 -1009
rect 281 -1040 320 -1030
rect 350 -1067 367 -977
rect 479 -1067 500 -867
rect 651 -884 668 -867
rect 805 -884 822 -867
rect 593 -892 634 -884
rect 593 -913 603 -892
rect 624 -913 634 -892
rect 651 -902 822 -884
rect 593 -922 634 -913
rect 805 -920 822 -902
rect 877 -920 915 -910
rect 805 -938 889 -920
rect 907 -938 915 -920
rect 665 -949 706 -940
rect 665 -970 677 -949
rect 698 -970 706 -949
rect 665 -978 706 -970
rect 736 -1009 775 -1002
rect 736 -1030 746 -1009
rect 767 -1030 775 -1009
rect 736 -1040 775 -1030
rect -619 -1079 -575 -1067
rect -619 -1120 -610 -1079
rect -588 -1120 -575 -1079
rect -619 -1132 -575 -1120
rect -556 -1079 -511 -1067
rect -556 -1120 -543 -1079
rect -521 -1120 -511 -1079
rect -556 -1132 -511 -1120
rect -482 -1079 -438 -1067
rect -482 -1120 -473 -1079
rect -451 -1120 -438 -1079
rect -482 -1132 -438 -1120
rect -419 -1079 -374 -1067
rect -419 -1120 -406 -1079
rect -384 -1120 -374 -1079
rect -419 -1132 -374 -1120
rect -336 -1080 -290 -1067
rect -336 -1121 -321 -1080
rect -299 -1121 -290 -1080
rect -336 -1132 -290 -1121
rect -131 -1078 -85 -1067
rect -131 -1119 -120 -1078
rect -98 -1119 -85 -1078
rect -131 -1132 -85 -1119
rect -50 -1079 -5 -1067
rect -50 -1120 -40 -1079
rect -18 -1120 -5 -1079
rect -50 -1132 -5 -1120
rect 14 -1079 59 -1067
rect 14 -1120 27 -1079
rect 49 -1120 59 -1079
rect 14 -1132 59 -1120
rect 116 -1080 162 -1067
rect 116 -1121 131 -1080
rect 153 -1121 162 -1080
rect 116 -1132 162 -1121
rect 321 -1078 367 -1067
rect 321 -1119 332 -1078
rect 354 -1119 367 -1078
rect 321 -1132 367 -1119
rect 402 -1079 447 -1067
rect 402 -1120 412 -1079
rect 434 -1120 447 -1079
rect 402 -1132 447 -1120
rect 466 -1079 511 -1067
rect 466 -1120 479 -1079
rect 501 -1120 511 -1079
rect 466 -1132 511 -1120
rect 571 -1080 617 -1067
rect 736 -1079 755 -1040
rect 805 -1067 822 -938
rect 877 -946 915 -938
rect 934 -1067 955 -867
rect 1101 -884 1118 -867
rect 1255 -884 1272 -867
rect 1043 -892 1084 -884
rect 1043 -913 1053 -892
rect 1074 -913 1084 -892
rect 1101 -902 1272 -884
rect 1043 -922 1084 -913
rect 1115 -949 1156 -940
rect 1115 -970 1127 -949
rect 1148 -970 1156 -949
rect 1115 -978 1156 -970
rect 1255 -961 1272 -902
rect 1320 -958 1357 -950
rect 1320 -961 1330 -958
rect 1255 -976 1330 -961
rect 1348 -976 1357 -958
rect 1126 -1046 1147 -978
rect 1255 -980 1357 -976
rect 1186 -1009 1225 -1002
rect 1186 -1030 1196 -1009
rect 1217 -1030 1225 -1009
rect 1186 -1040 1225 -1030
rect 1121 -1055 1155 -1046
rect 571 -1121 586 -1080
rect 608 -1121 617 -1080
rect 725 -1087 755 -1079
rect 725 -1104 733 -1087
rect 750 -1104 755 -1087
rect 725 -1110 755 -1104
rect 776 -1078 822 -1067
rect 571 -1132 617 -1121
rect 776 -1119 787 -1078
rect 809 -1119 822 -1078
rect 776 -1132 822 -1119
rect 857 -1079 902 -1067
rect 857 -1120 867 -1079
rect 889 -1120 902 -1079
rect 857 -1132 902 -1120
rect 921 -1079 966 -1067
rect 921 -1120 934 -1079
rect 956 -1120 966 -1079
rect 921 -1132 966 -1120
rect 1021 -1080 1067 -1067
rect 1021 -1121 1036 -1080
rect 1058 -1121 1067 -1080
rect 1121 -1072 1131 -1055
rect 1148 -1072 1155 -1055
rect 1255 -1067 1272 -980
rect 1320 -986 1357 -980
rect 1384 -1067 1405 -867
rect 1121 -1082 1155 -1072
rect 1226 -1078 1272 -1067
rect 1021 -1132 1067 -1121
rect 1226 -1119 1237 -1078
rect 1259 -1119 1272 -1078
rect 1226 -1132 1272 -1119
rect 1307 -1079 1352 -1067
rect 1307 -1120 1317 -1079
rect 1339 -1120 1352 -1079
rect 1307 -1132 1352 -1120
rect 1371 -1079 1416 -1067
rect 1371 -1120 1384 -1079
rect 1406 -1120 1416 -1079
rect 1371 -1132 1416 -1120
rect -611 -1181 -589 -1132
rect -474 -1181 -452 -1132
rect -334 -1181 -313 -1132
rect -41 -1181 -19 -1132
rect 118 -1181 139 -1132
rect 411 -1181 433 -1132
rect 573 -1181 594 -1132
rect 866 -1181 888 -1132
rect 1023 -1181 1044 -1132
rect 1316 -1181 1338 -1132
rect -619 -1186 1437 -1181
rect -619 -1187 -290 -1186
rect -619 -1208 -608 -1187
rect -587 -1208 -575 -1187
rect -554 -1208 -534 -1187
rect -513 -1208 -471 -1187
rect -450 -1208 -438 -1187
rect -417 -1208 -397 -1187
rect -376 -1208 -332 -1187
rect -311 -1207 -290 -1187
rect -269 -1187 -203 -1186
rect -269 -1207 -247 -1187
rect -311 -1208 -247 -1207
rect -226 -1207 -203 -1187
rect -182 -1207 -159 -1186
rect -138 -1187 162 -1186
rect -138 -1207 -119 -1187
rect -226 -1208 -119 -1207
rect -98 -1208 -75 -1187
rect -54 -1208 -38 -1187
rect -17 -1208 -5 -1187
rect 16 -1208 36 -1187
rect 57 -1208 120 -1187
rect 141 -1207 162 -1187
rect 183 -1187 249 -1186
rect 183 -1207 205 -1187
rect 141 -1208 205 -1207
rect 226 -1207 249 -1187
rect 270 -1207 293 -1186
rect 314 -1187 617 -1186
rect 314 -1207 333 -1187
rect 226 -1208 333 -1207
rect 354 -1208 377 -1187
rect 398 -1208 414 -1187
rect 435 -1208 447 -1187
rect 468 -1208 488 -1187
rect 509 -1208 575 -1187
rect 596 -1207 617 -1187
rect 638 -1187 704 -1186
rect 638 -1207 660 -1187
rect 596 -1208 660 -1207
rect 681 -1207 704 -1187
rect 725 -1207 748 -1186
rect 769 -1187 1067 -1186
rect 769 -1207 788 -1187
rect 681 -1208 788 -1207
rect 809 -1208 832 -1187
rect 853 -1208 869 -1187
rect 890 -1208 902 -1187
rect 923 -1208 943 -1187
rect 964 -1208 1025 -1187
rect 1046 -1207 1067 -1187
rect 1088 -1187 1154 -1186
rect 1088 -1207 1110 -1187
rect 1046 -1208 1110 -1207
rect 1131 -1207 1154 -1187
rect 1175 -1207 1198 -1186
rect 1219 -1187 1437 -1186
rect 1219 -1207 1238 -1187
rect 1131 -1208 1238 -1207
rect 1259 -1208 1282 -1187
rect 1303 -1208 1319 -1187
rect 1340 -1208 1352 -1187
rect 1373 -1208 1393 -1187
rect 1414 -1208 1437 -1187
rect -619 -1214 1437 -1208
rect -619 -1216 573 -1214
rect 594 -1216 1023 -1214
rect 1044 -1216 1437 -1214
rect -490 -1255 1457 -1251
rect -490 -1257 -88 -1255
rect -490 -1278 -476 -1257
rect -455 -1278 -434 -1257
rect -413 -1258 -323 -1257
rect -413 -1278 -395 -1258
rect -490 -1279 -395 -1278
rect -374 -1278 -323 -1258
rect -302 -1278 -280 -1257
rect -259 -1258 -145 -1257
rect -259 -1278 -236 -1258
rect -374 -1279 -236 -1278
rect -215 -1279 -191 -1258
rect -170 -1278 -145 -1258
rect -124 -1276 -88 -1257
rect -67 -1257 366 -1255
rect -67 -1276 -39 -1257
rect -124 -1278 -39 -1276
rect -18 -1278 3 -1257
rect 24 -1258 131 -1257
rect 24 -1278 42 -1258
rect -170 -1279 42 -1278
rect 63 -1278 131 -1258
rect 152 -1278 174 -1257
rect 195 -1258 309 -1257
rect 195 -1278 218 -1258
rect 63 -1279 218 -1278
rect 239 -1279 263 -1258
rect 284 -1278 309 -1258
rect 330 -1276 366 -1257
rect 387 -1257 821 -1255
rect 387 -1276 415 -1257
rect 330 -1278 415 -1276
rect 436 -1278 457 -1257
rect 478 -1258 586 -1257
rect 478 -1278 496 -1258
rect 284 -1279 496 -1278
rect 517 -1278 586 -1258
rect 607 -1278 629 -1257
rect 650 -1258 764 -1257
rect 650 -1278 673 -1258
rect 517 -1279 673 -1278
rect 694 -1279 718 -1258
rect 739 -1278 764 -1258
rect 785 -1276 821 -1257
rect 842 -1257 1276 -1255
rect 842 -1276 870 -1257
rect 785 -1278 870 -1276
rect 891 -1278 912 -1257
rect 933 -1258 1041 -1257
rect 933 -1278 951 -1258
rect 739 -1279 951 -1278
rect 972 -1278 1041 -1258
rect 1062 -1278 1084 -1257
rect 1105 -1258 1219 -1257
rect 1105 -1278 1128 -1258
rect 972 -1279 1128 -1278
rect 1149 -1278 1219 -1258
rect 1240 -1276 1276 -1257
rect 1297 -1257 1457 -1255
rect 1297 -1276 1325 -1257
rect 1240 -1278 1325 -1276
rect 1346 -1278 1367 -1257
rect 1388 -1258 1457 -1257
rect 1388 -1278 1406 -1258
rect 1149 -1279 1406 -1278
rect 1427 -1279 1457 -1258
rect -490 -1286 1457 -1279
rect -476 -1355 -455 -1286
rect -415 -1310 -356 -1303
rect -415 -1328 -384 -1310
rect -364 -1328 -356 -1310
rect -415 -1338 -356 -1328
rect -415 -1355 -395 -1338
rect -326 -1355 -301 -1286
rect -247 -1309 -209 -1303
rect -247 -1329 -239 -1309
rect -217 -1329 -209 -1309
rect -247 -1338 -209 -1329
rect -192 -1355 -167 -1286
rect -39 -1355 -18 -1286
rect 128 -1355 153 -1286
rect 262 -1355 287 -1286
rect 415 -1355 436 -1286
rect 583 -1355 608 -1286
rect 717 -1355 742 -1286
rect 870 -1355 891 -1286
rect 1038 -1355 1063 -1286
rect 1172 -1355 1197 -1286
rect 1325 -1355 1346 -1286
rect -490 -1371 -446 -1355
rect -490 -1406 -477 -1371
rect -452 -1406 -446 -1371
rect -490 -1419 -446 -1406
rect -427 -1371 -382 -1355
rect -427 -1406 -415 -1371
rect -390 -1406 -382 -1371
rect -427 -1419 -382 -1406
rect -341 -1370 -294 -1355
rect -341 -1405 -328 -1370
rect -303 -1405 -294 -1370
rect -341 -1419 -294 -1405
rect -275 -1368 -225 -1355
rect -275 -1403 -262 -1368
rect -237 -1403 -225 -1368
rect -275 -1419 -225 -1403
rect -206 -1369 -154 -1355
rect -206 -1404 -193 -1369
rect -168 -1404 -154 -1369
rect -206 -1419 -154 -1404
rect -135 -1370 -88 -1355
rect -135 -1405 -125 -1370
rect -100 -1405 -88 -1370
rect -135 -1419 -88 -1405
rect -53 -1371 -9 -1355
rect -53 -1406 -40 -1371
rect -15 -1406 -9 -1371
rect -53 -1419 -9 -1406
rect 10 -1371 55 -1355
rect 10 -1406 22 -1371
rect 47 -1406 55 -1371
rect 10 -1419 55 -1406
rect 113 -1370 160 -1355
rect 113 -1405 126 -1370
rect 151 -1405 160 -1370
rect 113 -1419 160 -1405
rect 179 -1368 229 -1355
rect 179 -1403 192 -1368
rect 217 -1403 229 -1368
rect 179 -1419 229 -1403
rect 248 -1369 300 -1355
rect 248 -1404 261 -1369
rect 286 -1404 300 -1369
rect 248 -1419 300 -1404
rect 319 -1370 366 -1355
rect 319 -1405 329 -1370
rect 354 -1405 366 -1370
rect 319 -1419 366 -1405
rect 401 -1371 445 -1355
rect 401 -1406 414 -1371
rect 439 -1406 445 -1371
rect 401 -1419 445 -1406
rect 464 -1371 509 -1355
rect 464 -1406 476 -1371
rect 501 -1406 509 -1371
rect 464 -1419 509 -1406
rect 568 -1370 615 -1355
rect 568 -1405 581 -1370
rect 606 -1405 615 -1370
rect 568 -1419 615 -1405
rect 634 -1368 684 -1355
rect 634 -1403 647 -1368
rect 672 -1403 684 -1368
rect 634 -1419 684 -1403
rect 703 -1369 755 -1355
rect 703 -1404 716 -1369
rect 741 -1404 755 -1369
rect 703 -1419 755 -1404
rect 774 -1370 821 -1355
rect 774 -1405 784 -1370
rect 809 -1405 821 -1370
rect 774 -1419 821 -1405
rect 856 -1371 900 -1355
rect 856 -1406 869 -1371
rect 894 -1406 900 -1371
rect 856 -1419 900 -1406
rect 919 -1371 964 -1355
rect 919 -1406 931 -1371
rect 956 -1406 964 -1371
rect 919 -1419 964 -1406
rect 1023 -1370 1070 -1355
rect 1023 -1405 1036 -1370
rect 1061 -1405 1070 -1370
rect 1023 -1419 1070 -1405
rect 1089 -1368 1139 -1355
rect 1089 -1403 1102 -1368
rect 1127 -1403 1139 -1368
rect 1089 -1419 1139 -1403
rect 1158 -1369 1210 -1355
rect 1158 -1404 1171 -1369
rect 1196 -1404 1210 -1369
rect 1158 -1419 1210 -1404
rect 1229 -1370 1276 -1355
rect 1229 -1405 1239 -1370
rect 1264 -1405 1276 -1370
rect 1229 -1419 1276 -1405
rect 1311 -1371 1355 -1355
rect 1311 -1406 1324 -1371
rect 1349 -1406 1355 -1371
rect 1311 -1419 1355 -1406
rect 1374 -1371 1419 -1355
rect 1374 -1406 1386 -1371
rect 1411 -1406 1419 -1371
rect 1374 -1419 1419 -1406
rect -463 -1564 -431 -1555
rect -463 -1581 -454 -1564
rect -437 -1581 -431 -1564
rect -463 -1589 -431 -1581
rect -414 -1566 -393 -1419
rect -260 -1436 -243 -1419
rect -106 -1436 -89 -1419
rect -318 -1444 -277 -1436
rect -318 -1465 -308 -1444
rect -287 -1465 -277 -1444
rect -260 -1454 -89 -1436
rect -318 -1474 -277 -1465
rect -175 -1561 -136 -1554
rect -175 -1566 -165 -1561
rect -414 -1582 -165 -1566
rect -144 -1582 -136 -1561
rect -414 -1584 -136 -1582
rect -414 -1619 -393 -1584
rect -175 -1592 -136 -1584
rect -106 -1576 -89 -1454
rect -31 -1574 2 -1569
rect -31 -1576 -23 -1574
rect -106 -1591 -23 -1576
rect -6 -1591 2 -1574
rect -106 -1593 2 -1591
rect -106 -1619 -89 -1593
rect -31 -1599 2 -1593
rect 23 -1619 44 -1419
rect 194 -1436 211 -1419
rect 348 -1436 365 -1419
rect 136 -1444 177 -1436
rect 136 -1465 146 -1444
rect 167 -1465 177 -1444
rect 194 -1454 365 -1436
rect 136 -1474 177 -1465
rect 208 -1501 249 -1492
rect 208 -1522 220 -1501
rect 241 -1522 249 -1501
rect 208 -1530 249 -1522
rect 219 -1558 239 -1530
rect 200 -1568 242 -1558
rect 200 -1589 211 -1568
rect 233 -1589 242 -1568
rect 200 -1598 242 -1589
rect 279 -1561 318 -1554
rect 279 -1582 289 -1561
rect 310 -1582 318 -1561
rect 279 -1592 318 -1582
rect 348 -1566 365 -1454
rect 417 -1564 451 -1555
rect 417 -1566 425 -1564
rect 348 -1581 425 -1566
rect 443 -1581 451 -1564
rect 348 -1583 451 -1581
rect 348 -1619 365 -1583
rect 417 -1588 451 -1583
rect 477 -1619 498 -1419
rect 649 -1436 666 -1419
rect 803 -1436 820 -1419
rect 591 -1444 632 -1436
rect 591 -1465 601 -1444
rect 622 -1465 632 -1444
rect 649 -1454 820 -1436
rect 591 -1474 632 -1465
rect 663 -1501 704 -1492
rect 663 -1522 675 -1501
rect 696 -1522 704 -1501
rect 663 -1530 704 -1522
rect 730 -1563 773 -1554
rect 730 -1584 740 -1563
rect 765 -1584 773 -1563
rect 730 -1593 773 -1584
rect 803 -1569 820 -1454
rect 873 -1564 907 -1556
rect 873 -1569 882 -1564
rect 803 -1582 882 -1569
rect 900 -1582 907 -1564
rect 803 -1586 907 -1582
rect 803 -1619 820 -1586
rect 873 -1590 907 -1586
rect 932 -1619 953 -1419
rect 1104 -1436 1121 -1419
rect 1258 -1436 1275 -1419
rect 1046 -1444 1087 -1436
rect 1046 -1465 1056 -1444
rect 1077 -1465 1087 -1444
rect 1104 -1454 1275 -1436
rect 1046 -1474 1087 -1465
rect 1118 -1501 1159 -1492
rect 1118 -1522 1130 -1501
rect 1151 -1522 1159 -1501
rect 1118 -1530 1159 -1522
rect 1189 -1561 1228 -1554
rect 1189 -1582 1199 -1561
rect 1220 -1582 1228 -1561
rect 1189 -1592 1228 -1582
rect 1258 -1565 1275 -1454
rect 1326 -1565 1360 -1557
rect 1258 -1583 1335 -1565
rect 1353 -1583 1360 -1565
rect 1258 -1585 1360 -1583
rect 1258 -1619 1275 -1585
rect 1326 -1591 1360 -1585
rect 1387 -1619 1408 -1419
rect -490 -1631 -446 -1619
rect -490 -1672 -481 -1631
rect -459 -1672 -446 -1631
rect -490 -1684 -446 -1672
rect -427 -1631 -382 -1619
rect -427 -1672 -414 -1631
rect -392 -1672 -382 -1631
rect -427 -1684 -382 -1672
rect -340 -1632 -294 -1619
rect -340 -1673 -325 -1632
rect -303 -1673 -294 -1632
rect -340 -1684 -294 -1673
rect -135 -1630 -89 -1619
rect -135 -1671 -124 -1630
rect -102 -1671 -89 -1630
rect -135 -1684 -89 -1671
rect -54 -1631 -9 -1619
rect -54 -1672 -44 -1631
rect -22 -1672 -9 -1631
rect -54 -1684 -9 -1672
rect 10 -1631 55 -1619
rect 10 -1672 23 -1631
rect 45 -1672 55 -1631
rect 10 -1684 55 -1672
rect 114 -1632 160 -1619
rect 114 -1673 129 -1632
rect 151 -1673 160 -1632
rect 114 -1684 160 -1673
rect 319 -1630 365 -1619
rect 319 -1671 330 -1630
rect 352 -1671 365 -1630
rect 319 -1684 365 -1671
rect 400 -1631 445 -1619
rect 400 -1672 410 -1631
rect 432 -1672 445 -1631
rect 400 -1684 445 -1672
rect 464 -1631 509 -1619
rect 464 -1672 477 -1631
rect 499 -1672 509 -1631
rect 464 -1684 509 -1672
rect 569 -1632 615 -1619
rect 569 -1673 584 -1632
rect 606 -1673 615 -1632
rect 569 -1684 615 -1673
rect 774 -1630 820 -1619
rect 774 -1671 785 -1630
rect 807 -1671 820 -1630
rect 774 -1684 820 -1671
rect 855 -1631 900 -1619
rect 855 -1672 865 -1631
rect 887 -1672 900 -1631
rect 855 -1684 900 -1672
rect 919 -1631 964 -1619
rect 919 -1672 932 -1631
rect 954 -1672 964 -1631
rect 919 -1684 964 -1672
rect 1024 -1632 1070 -1619
rect 1024 -1673 1039 -1632
rect 1061 -1673 1070 -1632
rect 1024 -1684 1070 -1673
rect 1229 -1630 1275 -1619
rect 1229 -1671 1240 -1630
rect 1262 -1671 1275 -1630
rect 1229 -1684 1275 -1671
rect 1310 -1631 1355 -1619
rect 1310 -1672 1320 -1631
rect 1342 -1672 1355 -1631
rect 1310 -1684 1355 -1672
rect 1374 -1631 1419 -1619
rect 1374 -1672 1387 -1631
rect 1409 -1672 1419 -1631
rect 1374 -1684 1419 -1672
rect -482 -1733 -460 -1684
rect -338 -1733 -317 -1684
rect -45 -1733 -23 -1684
rect 116 -1733 137 -1684
rect 409 -1733 431 -1684
rect 571 -1733 592 -1684
rect 864 -1733 886 -1684
rect 1026 -1733 1047 -1684
rect 1319 -1733 1341 -1684
rect -490 -1738 1452 -1733
rect -490 -1739 -294 -1738
rect -490 -1760 -479 -1739
rect -458 -1760 -446 -1739
rect -425 -1760 -405 -1739
rect -384 -1760 -336 -1739
rect -315 -1759 -294 -1739
rect -273 -1739 -207 -1738
rect -273 -1759 -251 -1739
rect -315 -1760 -251 -1759
rect -230 -1759 -207 -1739
rect -186 -1759 -163 -1738
rect -142 -1739 160 -1738
rect -142 -1759 -123 -1739
rect -230 -1760 -123 -1759
rect -102 -1760 -79 -1739
rect -58 -1760 -42 -1739
rect -21 -1760 -9 -1739
rect 12 -1760 32 -1739
rect 53 -1760 118 -1739
rect 139 -1759 160 -1739
rect 181 -1739 247 -1738
rect 181 -1759 203 -1739
rect 139 -1760 203 -1759
rect 224 -1759 247 -1739
rect 268 -1759 291 -1738
rect 312 -1739 615 -1738
rect 312 -1759 331 -1739
rect 224 -1760 331 -1759
rect 352 -1760 375 -1739
rect 396 -1760 412 -1739
rect 433 -1760 445 -1739
rect 466 -1760 486 -1739
rect 507 -1760 573 -1739
rect 594 -1759 615 -1739
rect 636 -1739 702 -1738
rect 636 -1759 658 -1739
rect 594 -1760 658 -1759
rect 679 -1759 702 -1739
rect 723 -1759 746 -1738
rect 767 -1739 1070 -1738
rect 767 -1759 786 -1739
rect 679 -1760 786 -1759
rect 807 -1760 830 -1739
rect 851 -1760 867 -1739
rect 888 -1760 900 -1739
rect 921 -1760 941 -1739
rect 962 -1760 1028 -1739
rect 1049 -1759 1070 -1739
rect 1091 -1739 1157 -1738
rect 1091 -1759 1113 -1739
rect 1049 -1760 1113 -1759
rect 1134 -1759 1157 -1739
rect 1178 -1759 1201 -1738
rect 1222 -1739 1452 -1738
rect 1222 -1759 1241 -1739
rect 1134 -1760 1241 -1759
rect 1262 -1760 1285 -1739
rect 1306 -1760 1322 -1739
rect 1343 -1760 1355 -1739
rect 1376 -1760 1396 -1739
rect 1417 -1760 1452 -1739
rect -490 -1766 1452 -1760
rect -490 -1768 -338 -1766
rect -317 -1768 116 -1766
rect 137 -1768 571 -1766
rect 592 -1768 1026 -1766
rect 1047 -1768 1452 -1766
<< viali >>
rect -605 -726 -584 -705
rect -468 -726 -447 -705
rect -319 -726 -298 -705
rect -187 -727 -166 -706
rect -35 -726 -14 -705
rect 133 -726 154 -705
rect 265 -727 286 -706
rect 417 -726 438 -705
rect 588 -726 609 -705
rect 720 -727 741 -706
rect 872 -726 893 -705
rect 1038 -726 1059 -705
rect 1170 -727 1191 -706
rect 1322 -726 1343 -705
rect -530 -912 -511 -895
rect -638 -982 -621 -965
rect -304 -913 -283 -892
rect -230 -970 -209 -949
rect -456 -1011 -431 -989
rect -161 -1030 -140 -1009
rect 148 -913 169 -892
rect 222 -970 243 -949
rect 291 -1030 312 -1009
rect 603 -913 624 -892
rect 677 -970 698 -949
rect 1053 -913 1074 -892
rect 1127 -970 1148 -949
rect 1196 -1030 1217 -1009
rect 733 -1104 750 -1087
rect 1131 -1072 1148 -1055
rect -608 -1208 -587 -1187
rect -471 -1208 -450 -1187
rect -332 -1208 -311 -1187
rect -38 -1208 -17 -1187
rect 120 -1208 141 -1187
rect 414 -1208 435 -1187
rect 575 -1208 596 -1187
rect 869 -1208 890 -1187
rect 1025 -1208 1046 -1187
rect 1319 -1208 1340 -1187
rect -476 -1278 -455 -1257
rect -323 -1278 -302 -1257
rect -191 -1279 -170 -1258
rect -39 -1278 -18 -1257
rect 131 -1278 152 -1257
rect 263 -1279 284 -1258
rect 415 -1278 436 -1257
rect 586 -1278 607 -1257
rect 718 -1279 739 -1258
rect 870 -1278 891 -1257
rect 1041 -1278 1062 -1257
rect 1325 -1278 1346 -1257
rect -384 -1328 -364 -1310
rect -239 -1329 -217 -1309
rect -454 -1581 -437 -1564
rect -308 -1465 -287 -1444
rect -165 -1582 -144 -1561
rect 146 -1465 167 -1444
rect 211 -1589 233 -1568
rect 289 -1582 310 -1561
rect 601 -1465 622 -1444
rect 675 -1522 696 -1501
rect 740 -1584 765 -1563
rect 1056 -1465 1077 -1444
rect 1130 -1522 1151 -1501
rect 1199 -1582 1220 -1561
rect -479 -1760 -458 -1739
rect -336 -1760 -315 -1739
rect -42 -1760 -21 -1739
rect 118 -1760 139 -1739
rect 412 -1760 433 -1739
rect 573 -1760 594 -1739
rect 867 -1760 888 -1739
rect 1028 -1760 1049 -1739
rect 1322 -1760 1343 -1739
<< metal1 >>
rect -619 -705 1437 -699
rect -619 -726 -605 -705
rect -584 -726 -468 -705
rect -447 -726 -319 -705
rect -298 -706 -35 -705
rect -298 -726 -187 -706
rect -619 -727 -187 -726
rect -166 -726 -35 -706
rect -14 -726 133 -705
rect 154 -706 417 -705
rect 154 -726 265 -706
rect -166 -727 265 -726
rect 286 -726 417 -706
rect 438 -726 588 -705
rect 609 -706 872 -705
rect 609 -726 720 -706
rect 286 -727 720 -726
rect 741 -726 872 -706
rect 893 -726 1038 -705
rect 1059 -706 1322 -705
rect 1059 -726 1170 -706
rect 741 -727 1170 -726
rect 1191 -726 1322 -706
rect 1343 -726 1437 -705
rect 1191 -727 1437 -726
rect -619 -734 1437 -727
rect -541 -895 -500 -885
rect -314 -892 -273 -884
rect -314 -895 -304 -892
rect -541 -912 -530 -895
rect -511 -912 -304 -895
rect -541 -913 -304 -912
rect -283 -895 -273 -892
rect 138 -892 179 -884
rect 138 -895 148 -892
rect -283 -913 148 -895
rect 169 -895 179 -892
rect 593 -892 634 -884
rect 593 -895 603 -892
rect 169 -913 603 -895
rect 624 -895 634 -892
rect 1043 -892 1084 -884
rect 1043 -895 1053 -892
rect 624 -913 1053 -895
rect 1074 -913 1084 -892
rect -541 -923 -500 -913
rect -314 -922 -273 -913
rect 138 -922 179 -913
rect 593 -922 634 -913
rect 1043 -922 1084 -913
rect -242 -944 -201 -940
rect -648 -965 -610 -957
rect -648 -982 -638 -965
rect -621 -982 -610 -965
rect -242 -974 -239 -944
rect -204 -953 -201 -944
rect 210 -945 251 -940
rect 210 -953 216 -945
rect -204 -967 216 -953
rect -204 -974 -201 -967
rect -242 -978 -201 -974
rect 210 -973 216 -967
rect 246 -973 251 -945
rect 210 -978 251 -973
rect 665 -949 706 -940
rect 665 -970 677 -949
rect 698 -953 706 -949
rect 1115 -949 1156 -940
rect 1115 -953 1127 -949
rect 698 -968 1127 -953
rect 698 -970 706 -968
rect 665 -978 706 -970
rect 1115 -970 1127 -968
rect 1148 -970 1156 -949
rect 1115 -978 1156 -970
rect -648 -990 -610 -982
rect -468 -984 -423 -980
rect -648 -1452 -633 -990
rect -468 -1017 -464 -984
rect -429 -1017 -423 -984
rect -171 -1009 -132 -1002
rect -171 -1017 -161 -1009
rect -468 -1022 -423 -1017
rect -381 -1030 -161 -1017
rect -140 -1030 -132 -1009
rect -381 -1033 -132 -1030
rect -619 -1187 -435 -1181
rect -619 -1208 -608 -1187
rect -587 -1208 -471 -1187
rect -450 -1208 -435 -1187
rect -619 -1216 -435 -1208
rect -490 -1257 -433 -1251
rect -490 -1278 -476 -1257
rect -455 -1278 -433 -1257
rect -490 -1286 -433 -1278
rect -381 -1303 -361 -1033
rect -171 -1040 -132 -1033
rect 281 -1009 320 -1002
rect 281 -1030 291 -1009
rect 312 -1010 320 -1009
rect 1186 -1009 1225 -1002
rect 1186 -1010 1196 -1009
rect 312 -1030 1196 -1010
rect 1217 -1015 1225 -1009
rect 1217 -1030 1280 -1015
rect 281 -1031 1280 -1030
rect 281 -1040 320 -1031
rect 1186 -1040 1225 -1031
rect -161 -1088 -142 -1040
rect 1121 -1055 1155 -1046
rect 1121 -1072 1131 -1055
rect 1148 -1072 1155 -1055
rect 725 -1087 755 -1079
rect 725 -1088 733 -1087
rect -161 -1104 733 -1088
rect 750 -1104 755 -1087
rect -161 -1109 755 -1104
rect 725 -1110 755 -1109
rect 1121 -1082 1155 -1072
rect -343 -1187 1079 -1181
rect -343 -1208 -332 -1187
rect -311 -1208 -38 -1187
rect -17 -1208 120 -1187
rect 141 -1208 414 -1187
rect 435 -1208 575 -1187
rect 596 -1208 869 -1187
rect 890 -1208 1025 -1187
rect 1046 -1208 1079 -1187
rect -343 -1216 1079 -1208
rect -336 -1257 1079 -1251
rect -336 -1278 -323 -1257
rect -302 -1258 -39 -1257
rect -302 -1278 -191 -1258
rect -336 -1279 -191 -1278
rect -170 -1278 -39 -1258
rect -18 -1278 131 -1257
rect 152 -1258 415 -1257
rect 152 -1278 263 -1258
rect -170 -1279 263 -1278
rect 284 -1278 415 -1258
rect 436 -1278 586 -1257
rect 607 -1258 870 -1257
rect 607 -1278 718 -1258
rect 284 -1279 718 -1278
rect 739 -1278 870 -1258
rect 891 -1278 1041 -1257
rect 1062 -1278 1079 -1257
rect 739 -1279 1079 -1278
rect -336 -1286 1079 -1279
rect -396 -1310 -356 -1303
rect -396 -1328 -384 -1310
rect -364 -1328 -356 -1310
rect -396 -1338 -356 -1328
rect -247 -1307 -206 -1303
rect -247 -1338 -239 -1307
rect -210 -1338 -206 -1307
rect -247 -1344 -206 -1338
rect -318 -1444 -277 -1436
rect -318 -1452 -308 -1444
rect -648 -1465 -308 -1452
rect -287 -1445 -277 -1444
rect 136 -1444 177 -1436
rect 136 -1445 146 -1444
rect -287 -1463 146 -1445
rect -287 -1465 -277 -1463
rect -648 -1466 -277 -1465
rect -318 -1474 -277 -1466
rect 136 -1465 146 -1463
rect 167 -1445 177 -1444
rect 591 -1444 632 -1436
rect 591 -1445 601 -1444
rect 167 -1463 601 -1445
rect 167 -1465 177 -1463
rect 136 -1474 177 -1465
rect 591 -1465 601 -1463
rect 622 -1445 632 -1444
rect 1046 -1444 1087 -1436
rect 1046 -1445 1056 -1444
rect 622 -1463 1056 -1445
rect 622 -1465 632 -1463
rect 591 -1474 632 -1465
rect 1046 -1465 1056 -1463
rect 1077 -1465 1087 -1444
rect 1046 -1474 1087 -1465
rect -534 -1496 -491 -1488
rect 1121 -1492 1147 -1082
rect -534 -1522 -528 -1496
rect -498 -1502 -491 -1496
rect 663 -1501 704 -1492
rect 663 -1502 675 -1501
rect -498 -1518 675 -1502
rect -498 -1522 -491 -1518
rect -534 -1527 -491 -1522
rect 663 -1522 675 -1518
rect 696 -1502 704 -1501
rect 1118 -1501 1159 -1492
rect 1118 -1502 1130 -1501
rect 696 -1518 1130 -1502
rect 696 -1522 704 -1518
rect 663 -1530 704 -1522
rect 1118 -1522 1130 -1518
rect 1151 -1522 1159 -1501
rect 1118 -1530 1159 -1522
rect -463 -1564 -431 -1555
rect -463 -1568 -454 -1564
rect -466 -1581 -454 -1568
rect -437 -1581 -431 -1564
rect -466 -1584 -431 -1581
rect -463 -1589 -431 -1584
rect -175 -1558 -136 -1554
rect -175 -1587 -169 -1558
rect -141 -1587 -136 -1558
rect -462 -1636 -439 -1589
rect -175 -1592 -136 -1587
rect 200 -1563 242 -1558
rect 200 -1592 207 -1563
rect 238 -1592 242 -1563
rect 279 -1561 318 -1554
rect 279 -1582 289 -1561
rect 310 -1582 318 -1561
rect 279 -1592 318 -1582
rect 730 -1560 773 -1554
rect 730 -1589 738 -1560
rect 768 -1589 773 -1560
rect 200 -1598 242 -1592
rect 290 -1636 308 -1592
rect 730 -1593 773 -1589
rect 1189 -1561 1228 -1554
rect 1189 -1582 1199 -1561
rect 1220 -1563 1228 -1561
rect 1255 -1563 1279 -1031
rect 1316 -1187 1437 -1181
rect 1316 -1208 1319 -1187
rect 1340 -1208 1437 -1187
rect 1316 -1216 1437 -1208
rect 1316 -1257 1457 -1251
rect 1316 -1278 1325 -1257
rect 1346 -1278 1457 -1257
rect 1316 -1286 1457 -1278
rect 1220 -1582 1279 -1563
rect 1189 -1584 1279 -1582
rect 1189 -1592 1228 -1584
rect 1189 -1636 1210 -1592
rect -462 -1656 1211 -1636
rect -490 -1739 1452 -1733
rect -490 -1760 -479 -1739
rect -458 -1760 -336 -1739
rect -315 -1760 -42 -1739
rect -21 -1760 118 -1739
rect 139 -1760 412 -1739
rect 433 -1760 573 -1739
rect 594 -1760 867 -1739
rect 888 -1760 1028 -1739
rect 1049 -1760 1322 -1739
rect 1343 -1760 1452 -1739
rect -490 -1768 1452 -1760
<< via1 >>
rect -239 -949 -204 -944
rect -239 -970 -230 -949
rect -230 -970 -209 -949
rect -209 -970 -204 -949
rect 216 -949 246 -945
rect -239 -974 -204 -970
rect 216 -970 222 -949
rect 222 -970 243 -949
rect 243 -970 246 -949
rect 216 -973 246 -970
rect -464 -989 -429 -984
rect -464 -1011 -456 -989
rect -456 -1011 -431 -989
rect -431 -1011 -429 -989
rect -464 -1017 -429 -1011
rect -239 -1309 -210 -1307
rect -239 -1329 -217 -1309
rect -217 -1329 -210 -1309
rect -239 -1338 -210 -1329
rect -528 -1522 -498 -1496
rect -169 -1561 -141 -1558
rect -169 -1582 -165 -1561
rect -165 -1582 -144 -1561
rect -144 -1582 -141 -1561
rect -169 -1587 -141 -1582
rect 207 -1568 238 -1563
rect 207 -1589 211 -1568
rect 211 -1589 233 -1568
rect 233 -1589 238 -1568
rect 207 -1592 238 -1589
rect 738 -1563 768 -1560
rect 738 -1584 740 -1563
rect 740 -1584 765 -1563
rect 765 -1584 768 -1563
rect 738 -1589 768 -1584
<< metal2 >>
rect -245 -944 -196 -938
rect -245 -974 -239 -944
rect -204 -974 -196 -944
rect -468 -984 -423 -980
rect -245 -982 -196 -974
rect 208 -945 251 -940
rect 208 -973 216 -945
rect 246 -973 251 -945
rect 208 -978 251 -973
rect -468 -993 -464 -984
rect -521 -1014 -464 -993
rect -521 -1488 -498 -1014
rect -468 -1017 -464 -1014
rect -429 -1017 -423 -984
rect -468 -1022 -423 -1017
rect -232 -1303 -213 -982
rect -247 -1307 -206 -1303
rect -247 -1338 -239 -1307
rect -210 -1338 -206 -1307
rect -247 -1344 -206 -1338
rect -534 -1496 -491 -1488
rect -534 -1522 -528 -1496
rect -498 -1522 -491 -1496
rect -534 -1527 -491 -1522
rect -175 -1558 -136 -1554
rect 208 -1558 231 -978
rect -175 -1587 -169 -1558
rect -141 -1587 -136 -1558
rect -175 -1592 -136 -1587
rect 200 -1563 242 -1558
rect 200 -1592 207 -1563
rect 238 -1592 242 -1563
rect -167 -1637 -147 -1592
rect 200 -1598 242 -1592
rect 730 -1560 773 -1554
rect 730 -1589 738 -1560
rect 768 -1589 773 -1560
rect 730 -1593 773 -1589
rect 743 -1637 759 -1593
rect -167 -1657 759 -1637
<< labels >>
flabel locali s -612 -732 -567 -704 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel locali s -487 -1285 -442 -1257 0 FreeSans 80 0 0 0 VDD
flabel locali s -615 -1214 -570 -1186 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel locali s -488 -1767 -443 -1739 0 FreeSans 80 0 0 0 GND
flabel poly s -598 -982 -553 -954 0 FreeSans 80 0 0 0 A
port 2 nsew
flabel poly s -456 -968 -411 -940 0 FreeSans 80 0 0 0 B
port 3 nsew
flabel poly s -462 -1551 -417 -1523 0 FreeSans 80 0 0 0 C
port 4 nsew
flabel locali s 21 -1037 53 -1002 0 FreeSans 80 0 0 0 O1
port 5 nsew
flabel locali s 479 -991 511 -956 0 FreeSans 80 0 0 0 O2
port 6 nsew
flabel locali s 930 -1006 962 -971 0 FreeSans 80 0 0 0 O3
port 7 nsew
flabel locali s 1378 -1027 1410 -992 0 FreeSans 80 0 0 0 O4
port 8 nsew
flabel locali s 20 -1599 52 -1564 0 FreeSans 80 0 0 0 O5
port 9 nsew
flabel locali s 472 -1591 504 -1556 0 FreeSans 80 0 0 0 O6
port 10 nsew
flabel locali s 924 -1592 956 -1557 0 FreeSans 80 0 0 0 O7
port 11 nsew
flabel locali s 1379 -1586 1411 -1551 0 FreeSans 80 0 0 0 O8
port 12 nsew
<< end >>
