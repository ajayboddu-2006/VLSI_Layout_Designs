magic

tech sky130A

timestamp 1738425198

<< nwell >>

rect -59 -13 2123 161

rect -57 -14 2123 -13

<< nmos >>

rect 1 -135 20 -83

rect 128 -135 147 -83

rect 256 -135 275 -83

rect 383 -135 402 -83

rect 511 -135 530 -83

rect 638 -135 657 -83

rect 766 -135 785 -83

rect 893 -135 912 -83

rect 1021 -135 1040 -83

rect 1152 -135 1171 -83

rect 1279 -135 1298 -83

rect 1407 -135 1426 -83

rect 1534 -135 1553 -83

rect 1662 -135 1681 -83

rect 1789 -135 1808 -83

rect 1917 -135 1936 -83

rect 2044 -135 2063 -83

<< pmos >>

rect 1 7 20 58

rect 128 7 147 58

rect 256 7 275 58

rect 383 7 402 58

rect 511 7 530 58

rect 638 7 657 58

rect 766 7 785 58

rect 893 7 912 58

rect 1021 7 1040 58

rect 1152 7 1171 58

rect 1279 7 1298 58

rect 1407 7 1426 58

rect 1534 7 1553 58

rect 1662 7 1681 58

rect 1789 7 1808 58

rect 1917 7 1936 58

rect 2044 7 2063 58

<< ndiff >>

rect -39 -90 1 -83

rect -39 -128 -31 -90

rect -9 -128 1 -90

rect -39 -135 1 -128

rect 20 -90 60 -83

rect 20 -128 30 -90

rect 52 -128 60 -90

rect 20 -135 60 -128

rect 88 -90 128 -83

rect 88 -128 96 -90

rect 118 -128 128 -90

rect 88 -135 128 -128

rect 147 -90 187 -83

rect 147 -128 157 -90

rect 179 -128 187 -90

rect 147 -135 187 -128

rect 216 -90 256 -83

rect 216 -128 224 -90

rect 246 -128 256 -90

rect 216 -135 256 -128

rect 275 -90 315 -83

rect 275 -128 285 -90

rect 307 -128 315 -90

rect 275 -135 315 -128

rect 343 -90 383 -83

rect 343 -128 351 -90

rect 373 -128 383 -90

rect 343 -135 383 -128

rect 402 -90 442 -83

rect 402 -128 412 -90

rect 434 -128 442 -90

rect 402 -135 442 -128

rect 471 -90 511 -83

rect 471 -128 479 -90

rect 501 -128 511 -90

rect 471 -135 511 -128

rect 530 -90 570 -83

rect 530 -128 540 -90

rect 562 -128 570 -90

rect 530 -135 570 -128

rect 598 -90 638 -83

rect 598 -128 606 -90

rect 628 -128 638 -90

rect 598 -135 638 -128

rect 657 -90 697 -83

rect 657 -128 667 -90

rect 689 -128 697 -90

rect 657 -135 697 -128

rect 726 -90 766 -83

rect 726 -128 734 -90

rect 756 -128 766 -90

rect 726 -135 766 -128

rect 785 -90 825 -83

rect 785 -128 795 -90

rect 817 -128 825 -90

rect 785 -135 825 -128

rect 853 -90 893 -83

rect 853 -128 861 -90

rect 883 -128 893 -90

rect 853 -135 893 -128

rect 912 -90 952 -83

rect 912 -128 922 -90

rect 944 -128 952 -90

rect 912 -135 952 -128

rect 981 -90 1021 -83

rect 981 -128 989 -90

rect 1011 -128 1021 -90

rect 981 -135 1021 -128

rect 1040 -90 1080 -83

rect 1040 -128 1050 -90

rect 1072 -128 1080 -90

rect 1040 -135 1080 -128

rect 1112 -90 1152 -83

rect 1112 -128 1120 -90

rect 1142 -128 1152 -90

rect 1112 -135 1152 -128

rect 1171 -90 1211 -83

rect 1171 -128 1181 -90

rect 1203 -128 1211 -90

rect 1171 -135 1211 -128

rect 1239 -90 1279 -83

rect 1239 -128 1247 -90

rect 1269 -128 1279 -90

rect 1239 -135 1279 -128

rect 1298 -90 1338 -83

rect 1298 -128 1308 -90

rect 1330 -128 1338 -90

rect 1298 -135 1338 -128

rect 1367 -90 1407 -83

rect 1367 -128 1375 -90

rect 1397 -128 1407 -90

rect 1367 -135 1407 -128

rect 1426 -90 1466 -83

rect 1426 -128 1436 -90

rect 1458 -128 1466 -90

rect 1426 -135 1466 -128

rect 1494 -90 1534 -83

rect 1494 -128 1502 -90

rect 1524 -128 1534 -90

rect 1494 -135 1534 -128

rect 1553 -90 1593 -83

rect 1553 -128 1563 -90

rect 1585 -128 1593 -90

rect 1553 -135 1593 -128

rect 1622 -90 1662 -83

rect 1622 -128 1630 -90

rect 1652 -128 1662 -90

rect 1622 -135 1662 -128

rect 1681 -90 1721 -83

rect 1681 -128 1691 -90

rect 1713 -128 1721 -90

rect 1681 -135 1721 -128

rect 1749 -90 1789 -83

rect 1749 -128 1757 -90

rect 1779 -128 1789 -90

rect 1749 -135 1789 -128

rect 1808 -90 1848 -83

rect 1808 -128 1818 -90

rect 1840 -128 1848 -90

rect 1808 -135 1848 -128

rect 1877 -90 1917 -83

rect 1877 -128 1885 -90

rect 1907 -128 1917 -90

rect 1877 -135 1917 -128

rect 1936 -90 1976 -83

rect 1936 -128 1946 -90

rect 1968 -128 1976 -90

rect 1936 -135 1976 -128

rect 2004 -90 2044 -83

rect 2004 -128 2012 -90

rect 2034 -128 2044 -90

rect 2004 -135 2044 -128

rect 2063 -90 2103 -83

rect 2063 -128 2073 -90

rect 2095 -128 2103 -90

rect 2063 -135 2103 -128

<< pdiff >>

rect -40 50 1 58

rect -40 15 -30 50

rect -6 15 1 50

rect -40 7 1 15

rect 20 50 61 58

rect 20 15 30 50

rect 54 15 61 50

rect 20 7 61 15

rect 88 50 128 58

rect 88 15 97 50

rect 121 15 128 50

rect 88 7 128 15

rect 147 50 188 58

rect 147 15 157 50

rect 181 15 188 50

rect 147 7 188 15

rect 215 50 256 58

rect 215 15 225 50

rect 249 15 256 50

rect 215 7 256 15

rect 275 50 316 58

rect 275 15 285 50

rect 309 15 316 50

rect 275 7 316 15

rect 343 50 383 58

rect 343 15 352 50

rect 376 15 383 50

rect 343 7 383 15

rect 402 50 443 58

rect 402 15 412 50

rect 436 15 443 50

rect 402 7 443 15

rect 470 50 511 58

rect 470 15 480 50

rect 504 15 511 50

rect 470 7 511 15

rect 530 50 571 58

rect 530 15 540 50

rect 564 15 571 50

rect 530 7 571 15

rect 598 50 638 58

rect 598 15 607 50

rect 631 15 638 50

rect 598 7 638 15

rect 657 50 698 58

rect 657 15 667 50

rect 691 15 698 50

rect 657 7 698 15

rect 725 50 766 58

rect 725 15 735 50

rect 759 15 766 50

rect 725 7 766 15

rect 785 50 826 58

rect 785 15 795 50

rect 819 15 826 50

rect 785 7 826 15

rect 853 50 893 58

rect 853 15 862 50

rect 886 15 893 50

rect 853 7 893 15

rect 912 50 953 58

rect 912 15 922 50

rect 946 15 953 50

rect 912 7 953 15

rect 980 50 1021 58

rect 980 15 990 50

rect 1014 15 1021 50

rect 980 7 1021 15

rect 1040 50 1081 58

rect 1040 15 1050 50

rect 1074 15 1081 50

rect 1040 7 1081 15

rect 1111 50 1152 58

rect 1111 15 1121 50

rect 1145 15 1152 50

rect 1111 7 1152 15

rect 1171 50 1212 58

rect 1171 15 1181 50

rect 1205 15 1212 50

rect 1171 7 1212 15

rect 1239 50 1279 58

rect 1239 15 1248 50

rect 1272 15 1279 50

rect 1239 7 1279 15

rect 1298 50 1339 58

rect 1298 15 1308 50

rect 1332 15 1339 50

rect 1298 7 1339 15

rect 1366 50 1407 58

rect 1366 15 1376 50

rect 1400 15 1407 50

rect 1366 7 1407 15

rect 1426 50 1467 58

rect 1426 15 1436 50

rect 1460 15 1467 50

rect 1426 7 1467 15

rect 1494 50 1534 58

rect 1494 15 1503 50

rect 1527 15 1534 50

rect 1494 7 1534 15

rect 1553 50 1594 58

rect 1553 15 1563 50

rect 1587 15 1594 50

rect 1553 7 1594 15

rect 1621 50 1662 58

rect 1621 15 1631 50

rect 1655 15 1662 50

rect 1621 7 1662 15

rect 1681 50 1722 58

rect 1681 15 1691 50

rect 1715 15 1722 50

rect 1681 7 1722 15

rect 1749 50 1789 58

rect 1749 15 1758 50

rect 1782 15 1789 50

rect 1749 7 1789 15

rect 1808 50 1849 58

rect 1808 15 1818 50

rect 1842 15 1849 50

rect 1808 7 1849 15

rect 1876 50 1917 58

rect 1876 15 1886 50

rect 1910 15 1917 50

rect 1876 7 1917 15

rect 1936 50 1977 58

rect 1936 15 1946 50

rect 1970 15 1977 50

rect 1936 7 1977 15

rect 2004 50 2044 58

rect 2004 15 2013 50

rect 2037 15 2044 50

rect 2004 7 2044 15

rect 2063 50 2104 58

rect 2063 15 2073 50

rect 2097 15 2104 50

rect 2063 7 2104 15

<< ndiffc >>

rect -31 -128 -9 -90

rect 30 -128 52 -90

rect 96 -128 118 -90

rect 157 -128 179 -90

rect 224 -128 246 -90

rect 285 -128 307 -90

rect 351 -128 373 -90

rect 412 -128 434 -90

rect 479 -128 501 -90

rect 540 -128 562 -90

rect 606 -128 628 -90

rect 667 -128 689 -90

rect 734 -128 756 -90

rect 795 -128 817 -90

rect 861 -128 883 -90

rect 922 -128 944 -90

rect 989 -128 1011 -90

rect 1050 -128 1072 -90

rect 1120 -128 1142 -90

rect 1181 -128 1203 -90

rect 1247 -128 1269 -90

rect 1308 -128 1330 -90

rect 1375 -128 1397 -90

rect 1436 -128 1458 -90

rect 1502 -128 1524 -90

rect 1563 -128 1585 -90

rect 1630 -128 1652 -90

rect 1691 -128 1713 -90

rect 1757 -128 1779 -90

rect 1818 -128 1840 -90

rect 1885 -128 1907 -90

rect 1946 -128 1968 -90

rect 2012 -128 2034 -90

rect 2073 -128 2095 -90

<< pdiffc >>

rect -30 15 -6 50

rect 30 15 54 50

rect 97 15 121 50

rect 157 15 181 50

rect 225 15 249 50

rect 285 15 309 50

rect 352 15 376 50

rect 412 15 436 50

rect 480 15 504 50

rect 540 15 564 50

rect 607 15 631 50

rect 667 15 691 50

rect 735 15 759 50

rect 795 15 819 50

rect 862 15 886 50

rect 922 15 946 50

rect 990 15 1014 50

rect 1050 15 1074 50

rect 1121 15 1145 50

rect 1181 15 1205 50

rect 1248 15 1272 50

rect 1308 15 1332 50

rect 1376 15 1400 50

rect 1436 15 1460 50

rect 1503 15 1527 50

rect 1563 15 1587 50

rect 1631 15 1655 50

rect 1691 15 1715 50

rect 1758 15 1782 50

rect 1818 15 1842 50

rect 1886 15 1910 50

rect 1946 15 1970 50

rect 2013 15 2037 50

rect 2073 15 2097 50

<< psubdiff >>

rect -58 -195 2122 -190

rect -58 -197 66 -195

rect -58 -217 6 -197

rect 26 -215 66 -197

rect 86 -215 134 -195

rect 154 -215 186 -195

rect 206 -197 579 -195

rect 206 -198 314 -197

rect 206 -215 268 -198

rect 26 -217 268 -215

rect -58 -218 268 -217

rect 288 -217 314 -198

rect 334 -217 395 -197

rect 415 -217 442 -197

rect 462 -217 527 -197

rect 547 -215 579 -197

rect 596 -215 644 -195

rect 664 -215 696 -195

rect 716 -197 1217 -195

rect 716 -198 824 -197

rect 716 -215 778 -198

rect 547 -217 778 -215

rect 288 -218 778 -217

rect 798 -217 824 -198

rect 844 -217 905 -197

rect 925 -217 952 -197

rect 972 -217 1037 -197

rect 1057 -217 1157 -197

rect 1177 -215 1217 -197

rect 1237 -215 1285 -195

rect 1305 -215 1337 -195

rect 1357 -197 1730 -195

rect 1357 -198 1465 -197

rect 1357 -215 1419 -198

rect 1177 -217 1419 -215

rect 798 -218 1419 -217

rect 1439 -217 1465 -198

rect 1485 -217 1546 -197

rect 1566 -217 1593 -197

rect 1613 -217 1678 -197

rect 1698 -215 1730 -197

rect 1747 -215 1795 -195

rect 1815 -215 1847 -195

rect 1867 -196 2122 -195

rect 1867 -197 2088 -196

rect 1867 -198 1975 -197

rect 1867 -215 1929 -198

rect 1698 -217 1929 -215

rect 1439 -218 1929 -217

rect 1949 -217 1975 -198

rect 1995 -217 2051 -197

rect 2071 -216 2088 -197

rect 2108 -216 2122 -196

rect 2071 -217 2122 -216

rect 1949 -218 2122 -217

rect -58 -221 2122 -218

<< nsubdiff >>

rect -40 138 1084 142

rect -40 137 134 138

rect -40 136 50 137

rect -40 116 7 136

rect 27 117 50 136

rect 70 118 134 137

rect 154 137 441 138

rect 154 118 179 137

rect 70 117 179 118

rect 199 117 260 137

rect 280 117 307 137

rect 327 136 441 137

rect 327 117 391 136

rect 27 116 391 117

rect 411 118 441 136

rect 461 136 644 138

rect 461 135 566 136

rect 461 118 522 135

rect 411 116 522 118

rect -40 115 522 116

rect 542 116 566 135

rect 586 118 644 136

rect 664 137 951 138

rect 664 118 689 137

rect 586 117 689 118

rect 709 117 770 137

rect 790 117 817 137

rect 837 136 951 137

rect 837 117 901 136

rect 586 116 901 117

rect 921 118 951 136

rect 971 135 1084 138

rect 971 118 1032 135

rect 921 116 1032 118

rect 542 115 1032 116

rect 1052 115 1084 135

rect -40 111 1084 115

rect 1111 138 2091 142

rect 1111 137 1285 138

rect 1111 136 1201 137

rect 1111 116 1158 136

rect 1178 117 1201 136

rect 1221 118 1285 137

rect 1305 137 1592 138

rect 1305 118 1330 137

rect 1221 117 1330 118

rect 1350 117 1411 137

rect 1431 117 1458 137

rect 1478 136 1592 137

rect 1478 117 1542 136

rect 1178 116 1542 117

rect 1562 118 1592 136

rect 1612 136 1795 138

rect 1612 135 1717 136

rect 1612 118 1673 135

rect 1562 116 1673 118

rect 1111 115 1673 116

rect 1693 116 1717 135

rect 1737 118 1795 136

rect 1815 137 2091 138

rect 1815 118 1840 137

rect 1737 117 1840 118

rect 1860 117 1921 137

rect 1941 117 1968 137

rect 1988 136 2091 137

rect 1988 117 2052 136

rect 1737 116 2052 117

rect 2072 116 2091 136

rect 1693 115 2091 116

rect 1111 111 2091 115

<< psubdiffcont >>

rect 6 -217 26 -197

rect 66 -215 86 -195

rect 134 -215 154 -195

rect 186 -215 206 -195

rect 268 -218 288 -198

rect 314 -217 334 -197

rect 395 -217 415 -197

rect 442 -217 462 -197

rect 527 -217 547 -197

rect 579 -215 596 -195

rect 644 -215 664 -195

rect 696 -215 716 -195

rect 778 -218 798 -198

rect 824 -217 844 -197

rect 905 -217 925 -197

rect 952 -217 972 -197

rect 1037 -217 1057 -197

rect 1157 -217 1177 -197

rect 1217 -215 1237 -195

rect 1285 -215 1305 -195

rect 1337 -215 1357 -195

rect 1419 -218 1439 -198

rect 1465 -217 1485 -197

rect 1546 -217 1566 -197

rect 1593 -217 1613 -197

rect 1678 -217 1698 -197

rect 1730 -215 1747 -195

rect 1795 -215 1815 -195

rect 1847 -215 1867 -195

rect 1929 -218 1949 -198

rect 1975 -217 1995 -197

rect 2051 -217 2071 -197

rect 2088 -216 2108 -196

<< nsubdiffcont >>

rect 7 116 27 136

rect 50 117 70 137

rect 134 118 154 138

rect 179 117 199 137

rect 260 117 280 137

rect 307 117 327 137

rect 391 116 411 136

rect 441 118 461 138

rect 522 115 542 135

rect 566 116 586 136

rect 644 118 664 138

rect 689 117 709 137

rect 770 117 790 137

rect 817 117 837 137

rect 901 116 921 136

rect 951 118 971 138

rect 1032 115 1052 135

rect 1158 116 1178 136

rect 1201 117 1221 137

rect 1285 118 1305 138

rect 1330 117 1350 137

rect 1411 117 1431 137

rect 1458 117 1478 137

rect 1542 116 1562 136

rect 1592 118 1612 138

rect 1673 115 1693 135

rect 1717 116 1737 136

rect 1795 118 1815 138

rect 1840 117 1860 137

rect 1921 117 1941 137

rect 1968 117 1988 137

rect 2052 116 2072 136

<< poly >>

rect 1 58 20 95

rect 128 58 147 95

rect 256 58 275 95

rect 383 58 402 95

rect 511 58 530 95

rect 638 58 657 95

rect 766 58 785 95

rect 893 58 912 95

rect 1021 58 1040 95

rect 1152 58 1171 95

rect 1279 58 1298 95

rect 1407 58 1426 95

rect 1534 58 1553 95

rect 1662 58 1681 95

rect 1789 58 1808 95

rect 1917 58 1936 95

rect 2044 58 2063 95

rect 1 -28 20 7

rect 128 -28 147 7

rect 256 -28 275 7

rect 383 -28 402 7

rect 511 -28 530 7

rect 638 -28 657 7

rect 766 -28 785 7

rect 893 -28 912 7

rect 1021 -28 1040 7

rect 1152 -28 1171 7

rect 1279 -28 1298 7

rect 1407 -28 1426 7

rect 1534 -28 1553 7

rect 1662 -28 1681 7

rect 1789 -28 1808 7

rect 1917 -28 1936 7

rect 2044 -28 2063 7

rect -34 -33 20 -28

rect -34 -53 -26 -33

rect -6 -53 20 -33

rect -34 -59 20 -53

rect 93 -33 147 -28

rect 93 -53 101 -33

rect 121 -53 147 -33

rect 93 -59 147 -53

rect 221 -33 275 -28

rect 221 -53 229 -33

rect 249 -53 275 -33

rect 221 -59 275 -53

rect 348 -33 402 -28

rect 348 -53 356 -33

rect 376 -53 402 -33

rect 348 -59 402 -53

rect 476 -33 530 -28

rect 476 -53 484 -33

rect 504 -53 530 -33

rect 476 -59 530 -53

rect 603 -33 657 -28

rect 603 -53 611 -33

rect 631 -53 657 -33

rect 603 -59 657 -53

rect 731 -33 785 -28

rect 731 -53 739 -33

rect 759 -53 785 -33

rect 731 -59 785 -53

rect 858 -33 912 -28

rect 858 -53 866 -33

rect 886 -53 912 -33

rect 858 -59 912 -53

rect 986 -33 1040 -28

rect 986 -53 994 -33

rect 1014 -53 1040 -33

rect 986 -59 1040 -53

rect 1117 -33 1171 -28

rect 1117 -53 1125 -33

rect 1145 -53 1171 -33

rect 1117 -59 1171 -53

rect 1244 -33 1298 -28

rect 1244 -53 1252 -33

rect 1272 -53 1298 -33

rect 1244 -59 1298 -53

rect 1372 -33 1426 -28

rect 1372 -53 1380 -33

rect 1400 -53 1426 -33

rect 1372 -59 1426 -53

rect 1499 -33 1553 -28

rect 1499 -53 1507 -33

rect 1527 -53 1553 -33

rect 1499 -59 1553 -53

rect 1627 -33 1681 -28

rect 1627 -53 1635 -33

rect 1655 -53 1681 -33

rect 1627 -59 1681 -53

rect 1754 -33 1808 -28

rect 1754 -53 1762 -33

rect 1782 -53 1808 -33

rect 1754 -59 1808 -53

rect 1882 -33 1936 -28

rect 1882 -53 1890 -33

rect 1910 -53 1936 -33

rect 1882 -59 1936 -53

rect 2009 -33 2063 -28

rect 2009 -53 2017 -33

rect 2037 -53 2063 -33

rect 2009 -59 2063 -53

rect 1 -83 20 -59

rect 128 -83 147 -59

rect 256 -83 275 -59

rect 383 -83 402 -59

rect 511 -83 530 -59

rect 638 -83 657 -59

rect 766 -83 785 -59

rect 893 -83 912 -59

rect 1021 -83 1040 -59

rect 1152 -83 1171 -59

rect 1279 -83 1298 -59

rect 1407 -83 1426 -59

rect 1534 -83 1553 -59

rect 1662 -83 1681 -59

rect 1789 -83 1808 -59

rect 1917 -83 1936 -59

rect 2044 -83 2063 -59

rect 1 -176 20 -135

rect 128 -176 147 -135

rect 256 -176 275 -135

rect 383 -176 402 -135

rect 511 -176 530 -135

rect 638 -176 657 -135

rect 766 -176 785 -135

rect 893 -176 912 -135

rect 1021 -176 1040 -135

rect 1152 -176 1171 -135

rect 1279 -176 1298 -135

rect 1407 -176 1426 -135

rect 1534 -176 1553 -135

rect 1662 -176 1681 -135

rect 1789 -176 1808 -135

rect 1917 -176 1936 -135

rect 2044 -176 2063 -135

<< polycont >>

rect -26 -53 -6 -33

rect 101 -53 121 -33

rect 229 -53 249 -33

rect 356 -53 376 -33

rect 484 -53 504 -33

rect 611 -53 631 -33

rect 739 -53 759 -33

rect 866 -53 886 -33

rect 994 -53 1014 -33

rect 1125 -53 1145 -33

rect 1252 -53 1272 -33

rect 1380 -53 1400 -33

rect 1507 -53 1527 -33

rect 1635 -53 1655 -33

rect 1762 -53 1782 -33

rect 1890 -53 1910 -33

rect 2017 -53 2037 -33

<< locali >>

rect -60 138 2123 142

rect -60 137 98 138

rect -60 136 50 137

rect -60 116 -30 136

rect -10 116 7 136

rect 27 117 50 136

rect 70 118 98 137

rect 118 118 134 138

rect 154 137 441 138

rect 154 118 179 137

rect 70 117 179 118

rect 199 117 221 137

rect 241 117 260 137

rect 280 117 307 137

rect 327 136 441 137

rect 327 117 350 136

rect 27 116 350 117

rect 370 116 391 136

rect 411 118 441 136

rect 461 136 608 138

rect 461 118 481 136

rect 411 116 481 118

rect 501 135 566 136

rect 501 116 522 135

rect -60 115 522 116

rect 542 116 566 135

rect 586 118 608 136

rect 628 118 644 138

rect 664 137 951 138

rect 664 118 689 137

rect 586 117 689 118

rect 709 117 731 137

rect 751 117 770 137

rect 790 117 817 137

rect 837 136 951 137

rect 837 117 860 136

rect 586 116 860 117

rect 880 116 901 136

rect 921 118 951 136

rect 971 137 1249 138

rect 971 136 1201 137

rect 971 118 991 136

rect 921 116 991 118

rect 1011 135 1121 136

rect 1011 116 1032 135

rect 542 115 1032 116

rect 1052 116 1121 135

rect 1141 116 1158 136

rect 1178 117 1201 136

rect 1221 118 1249 137

rect 1269 118 1285 138

rect 1305 137 1592 138

rect 1305 118 1330 137

rect 1221 117 1330 118

rect 1350 117 1372 137

rect 1392 117 1411 137

rect 1431 117 1458 137

rect 1478 136 1592 137

rect 1478 117 1501 136

rect 1178 116 1501 117

rect 1521 116 1542 136

rect 1562 118 1592 136

rect 1612 136 1759 138

rect 1612 118 1632 136

rect 1562 116 1632 118

rect 1652 135 1717 136

rect 1652 116 1673 135

rect 1052 115 1673 116

rect 1693 116 1717 135

rect 1737 118 1759 136

rect 1779 118 1795 138

rect 1815 137 2123 138

rect 1815 118 1840 137

rect 1737 117 1840 118

rect 1860 117 1882 137

rect 1902 117 1921 137

rect 1941 117 1968 137

rect 1988 136 2123 137

rect 1988 117 2011 136

rect 1737 116 2011 117

rect 2031 116 2052 136

rect 2072 116 2123 136

rect 1693 115 2123 116

rect -60 111 2123 115

rect -29 58 -9 111

rect 98 58 118 111

rect 225 58 245 111

rect 352 58 372 111

rect 481 58 501 111

rect 608 58 628 111

rect 735 58 755 111

rect 862 58 882 111

rect 991 58 1011 111

rect 1122 58 1142 111

rect 1249 58 1269 111

rect 1376 58 1396 111

rect 1503 58 1523 111

rect 1632 58 1652 111

rect 1759 58 1779 111

rect 1886 58 1906 111

rect 2013 58 2033 111

rect -40 50 -1 58

rect -40 15 -30 50

rect -6 15 -1 50

rect -40 7 -1 15

rect 22 50 61 58

rect 22 15 30 50

rect 54 15 61 50

rect 22 7 61 15

rect 88 50 126 58

rect 88 15 97 50

rect 121 15 126 50

rect 88 7 126 15

rect 149 50 188 58

rect 149 15 157 50

rect 181 15 188 50

rect 149 7 188 15

rect 215 50 254 58

rect 215 15 225 50

rect 249 15 254 50

rect 215 7 254 15

rect 277 50 316 58

rect 277 15 285 50

rect 309 15 316 50

rect 277 7 316 15

rect 343 50 381 58

rect 343 15 352 50

rect 376 15 381 50

rect 343 7 381 15

rect 404 50 443 58

rect 404 15 412 50

rect 436 15 443 50

rect 404 7 443 15

rect 470 50 509 58

rect 470 15 480 50

rect 504 15 509 50

rect 470 7 509 15

rect 532 50 571 58

rect 532 15 540 50

rect 564 15 571 50

rect 532 7 571 15

rect 598 50 636 58

rect 598 15 607 50

rect 631 15 636 50

rect 598 7 636 15

rect 659 50 698 58

rect 659 15 667 50

rect 691 15 698 50

rect 659 7 698 15

rect 725 50 764 58

rect 725 15 735 50

rect 759 15 764 50

rect 725 7 764 15

rect 787 50 826 58

rect 787 15 795 50

rect 819 15 826 50

rect 787 7 826 15

rect 853 50 891 58

rect 853 15 862 50

rect 886 15 891 50

rect 853 7 891 15

rect 914 50 953 58

rect 914 15 922 50

rect 946 15 953 50

rect 914 7 953 15

rect 980 50 1019 58

rect 980 15 990 50

rect 1014 15 1019 50

rect 980 7 1019 15

rect 1042 50 1081 58

rect 1042 15 1050 50

rect 1074 15 1081 50

rect 1042 7 1081 15

rect 1111 50 1150 58

rect 1111 15 1121 50

rect 1145 15 1150 50

rect 1111 7 1150 15

rect 1173 50 1212 58

rect 1173 15 1181 50

rect 1205 15 1212 50

rect 1173 7 1212 15

rect 1239 50 1277 58

rect 1239 15 1248 50

rect 1272 15 1277 50

rect 1239 7 1277 15

rect 1300 50 1339 58

rect 1300 15 1308 50

rect 1332 15 1339 50

rect 1300 7 1339 15

rect 1366 50 1405 58

rect 1366 15 1376 50

rect 1400 15 1405 50

rect 1366 7 1405 15

rect 1428 50 1467 58

rect 1428 15 1436 50

rect 1460 15 1467 50

rect 1428 7 1467 15

rect 1494 50 1532 58

rect 1494 15 1503 50

rect 1527 15 1532 50

rect 1494 7 1532 15

rect 1555 50 1594 58

rect 1555 15 1563 50

rect 1587 15 1594 50

rect 1555 7 1594 15

rect 1621 50 1660 58

rect 1621 15 1631 50

rect 1655 15 1660 50

rect 1621 7 1660 15

rect 1683 50 1722 58

rect 1683 15 1691 50

rect 1715 15 1722 50

rect 1683 7 1722 15

rect 1749 50 1787 58

rect 1749 15 1758 50

rect 1782 15 1787 50

rect 1749 7 1787 15

rect 1810 50 1849 58

rect 1810 15 1818 50

rect 1842 15 1849 50

rect 1810 7 1849 15

rect 1876 50 1915 58

rect 1876 15 1886 50

rect 1910 15 1915 50

rect 1876 7 1915 15

rect 1938 50 1977 58

rect 1938 15 1946 50

rect 1970 15 1977 50

rect 1938 7 1977 15

rect 2004 50 2042 58

rect 2004 15 2013 50

rect 2037 15 2042 50

rect 2004 7 2042 15

rect 2065 50 2104 58

rect 2065 15 2073 50

rect 2097 15 2104 50

rect 2065 7 2104 15

rect -34 -33 2 -28

rect -34 -53 -26 -33

rect -6 -53 2 -33

rect -34 -59 2 -53

rect 41 -33 60 7

rect 93 -33 129 -28

rect 41 -51 101 -33

rect 41 -83 60 -51

rect 93 -53 101 -51

rect 121 -53 129 -33

rect 93 -59 129 -53

rect 168 -33 187 7

rect 221 -33 257 -28

rect 168 -51 229 -33

rect 168 -83 187 -51

rect 221 -53 229 -51

rect 249 -53 257 -33

rect 221 -59 257 -53

rect 296 -33 315 7

rect 348 -33 384 -28

rect 296 -51 356 -33

rect 296 -83 315 -51

rect 348 -53 356 -51

rect 376 -53 384 -33

rect 348 -59 384 -53

rect 423 -32 442 7

rect 476 -32 512 -28

rect 423 -33 512 -32

rect 423 -50 484 -33

rect 423 -83 442 -50

rect 476 -53 484 -50

rect 504 -53 512 -33

rect 476 -59 512 -53

rect 551 -33 570 7

rect 603 -33 639 -28

rect 551 -51 611 -33

rect 551 -83 570 -51

rect 603 -53 611 -51

rect 631 -53 639 -33

rect 603 -59 639 -53

rect 678 -33 697 7

rect 731 -33 767 -28

rect 678 -51 739 -33

rect 678 -83 697 -51

rect 731 -53 739 -51

rect 759 -53 767 -33

rect 731 -59 767 -53

rect 806 -33 825 7

rect 858 -33 894 -28

rect 806 -51 866 -33

rect 806 -83 825 -51

rect 858 -53 866 -51

rect 886 -53 894 -33

rect 858 -59 894 -53

rect 933 -32 952 7

rect 986 -32 1022 -28

rect 933 -33 1022 -32

rect 933 -50 994 -33

rect 933 -83 952 -50

rect 986 -53 994 -50

rect 1014 -53 1022 -33

rect 986 -59 1022 -53

rect 1061 -35 1080 7

rect 1117 -33 1153 -28

rect 1117 -35 1125 -33

rect 1061 -52 1125 -35

rect 1061 -83 1080 -52

rect 1117 -53 1125 -52

rect 1145 -53 1153 -33

rect 1117 -59 1153 -53

rect 1192 -33 1211 7

rect 1244 -33 1280 -28

rect 1192 -51 1252 -33

rect 1192 -83 1211 -51

rect 1244 -53 1252 -51

rect 1272 -53 1280 -33

rect 1244 -59 1280 -53

rect 1319 -33 1338 7

rect 1372 -33 1408 -28

rect 1319 -51 1380 -33

rect 1319 -83 1338 -51

rect 1372 -53 1380 -51

rect 1400 -53 1408 -33

rect 1372 -59 1408 -53

rect 1447 -33 1466 7

rect 1499 -33 1535 -28

rect 1447 -51 1507 -33

rect 1447 -83 1466 -51

rect 1499 -53 1507 -51

rect 1527 -53 1535 -33

rect 1499 -59 1535 -53

rect 1574 -32 1593 7

rect 1627 -32 1663 -28

rect 1574 -33 1663 -32

rect 1574 -50 1635 -33

rect 1574 -83 1593 -50

rect 1627 -53 1635 -50

rect 1655 -53 1663 -33

rect 1627 -59 1663 -53

rect 1702 -33 1721 7

rect 1754 -33 1790 -28

rect 1702 -51 1762 -33

rect 1702 -83 1721 -51

rect 1754 -53 1762 -51

rect 1782 -53 1790 -33

rect 1754 -59 1790 -53

rect 1829 -33 1848 7

rect 1882 -33 1918 -28

rect 1829 -51 1890 -33

rect 1829 -83 1848 -51

rect 1882 -53 1890 -51

rect 1910 -53 1918 -33

rect 1882 -59 1918 -53

rect 1957 -33 1976 7

rect 2084 -26 2103 7

rect 2009 -33 2045 -28

rect 1957 -51 2017 -33

rect 1957 -83 1976 -51

rect 2009 -53 2017 -51

rect 2037 -53 2045 -33

rect 2009 -59 2045 -53

rect 2084 -30 2120 -26

rect 2084 -50 2093 -30

rect 2113 -50 2120 -30

rect 2084 -57 2120 -50

rect 2084 -83 2103 -57

rect -39 -90 -1 -83

rect -39 -128 -31 -90

rect -9 -128 -1 -90

rect -39 -135 -1 -128

rect 22 -90 60 -83

rect 22 -128 30 -90

rect 52 -128 60 -90

rect 22 -135 60 -128

rect 88 -90 126 -83

rect 88 -128 96 -90

rect 118 -128 126 -90

rect 88 -135 126 -128

rect 149 -90 187 -83

rect 149 -128 157 -90

rect 179 -128 187 -90

rect 149 -135 187 -128

rect 216 -90 254 -83

rect 216 -128 224 -90

rect 246 -128 254 -90

rect 216 -135 254 -128

rect 277 -90 315 -83

rect 277 -128 285 -90

rect 307 -128 315 -90

rect 277 -135 315 -128

rect 343 -90 381 -83

rect 343 -128 351 -90

rect 373 -128 381 -90

rect 343 -135 381 -128

rect 404 -90 442 -83

rect 404 -128 412 -90

rect 434 -128 442 -90

rect 404 -135 442 -128

rect 471 -90 509 -83

rect 471 -128 479 -90

rect 501 -128 509 -90

rect 471 -135 509 -128

rect 532 -90 570 -83

rect 532 -128 540 -90

rect 562 -128 570 -90

rect 532 -135 570 -128

rect 598 -90 636 -83

rect 598 -128 606 -90

rect 628 -128 636 -90

rect 598 -135 636 -128

rect 659 -90 697 -83

rect 659 -128 667 -90

rect 689 -128 697 -90

rect 659 -135 697 -128

rect 726 -90 764 -83

rect 726 -128 734 -90

rect 756 -128 764 -90

rect 726 -135 764 -128

rect 787 -90 825 -83

rect 787 -128 795 -90

rect 817 -128 825 -90

rect 787 -135 825 -128

rect 853 -90 891 -83

rect 853 -128 861 -90

rect 883 -128 891 -90

rect 853 -135 891 -128

rect 914 -90 952 -83

rect 914 -128 922 -90

rect 944 -128 952 -90

rect 914 -135 952 -128

rect 981 -90 1019 -83

rect 981 -128 989 -90

rect 1011 -128 1019 -90

rect 981 -135 1019 -128

rect 1042 -90 1080 -83

rect 1042 -128 1050 -90

rect 1072 -128 1080 -90

rect 1042 -135 1080 -128

rect 1112 -90 1150 -83

rect 1112 -128 1120 -90

rect 1142 -128 1150 -90

rect 1112 -135 1150 -128

rect 1173 -90 1211 -83

rect 1173 -128 1181 -90

rect 1203 -128 1211 -90

rect 1173 -135 1211 -128

rect 1239 -90 1277 -83

rect 1239 -128 1247 -90

rect 1269 -128 1277 -90

rect 1239 -135 1277 -128

rect 1300 -90 1338 -83

rect 1300 -128 1308 -90

rect 1330 -128 1338 -90

rect 1300 -135 1338 -128

rect 1367 -90 1405 -83

rect 1367 -128 1375 -90

rect 1397 -128 1405 -90

rect 1367 -135 1405 -128

rect 1428 -90 1466 -83

rect 1428 -128 1436 -90

rect 1458 -128 1466 -90

rect 1428 -135 1466 -128

rect 1494 -90 1532 -83

rect 1494 -128 1502 -90

rect 1524 -128 1532 -90

rect 1494 -135 1532 -128

rect 1555 -90 1593 -83

rect 1555 -128 1563 -90

rect 1585 -128 1593 -90

rect 1555 -135 1593 -128

rect 1622 -90 1660 -83

rect 1622 -128 1630 -90

rect 1652 -128 1660 -90

rect 1622 -135 1660 -128

rect 1683 -90 1721 -83

rect 1683 -128 1691 -90

rect 1713 -128 1721 -90

rect 1683 -135 1721 -128

rect 1749 -90 1787 -83

rect 1749 -128 1757 -90

rect 1779 -128 1787 -90

rect 1749 -135 1787 -128

rect 1810 -90 1848 -83

rect 1810 -128 1818 -90

rect 1840 -128 1848 -90

rect 1810 -135 1848 -128

rect 1877 -90 1915 -83

rect 1877 -128 1885 -90

rect 1907 -128 1915 -90

rect 1877 -135 1915 -128

rect 1938 -90 1976 -83

rect 1938 -128 1946 -90

rect 1968 -128 1976 -90

rect 1938 -135 1976 -128

rect 2004 -90 2042 -83

rect 2004 -128 2012 -90

rect 2034 -128 2042 -90

rect 2004 -135 2042 -128

rect 2065 -90 2103 -83

rect 2065 -128 2073 -90

rect 2095 -128 2103 -90

rect 2065 -135 2103 -128

rect -31 -190 -11 -135

rect 97 -190 117 -135

rect 225 -190 245 -135

rect 351 -190 374 -135

rect 478 -190 500 -135

rect 607 -190 627 -135

rect 735 -190 755 -135

rect 861 -190 884 -135

rect 988 -190 1010 -135

rect 1120 -190 1140 -135

rect 1248 -190 1268 -135

rect 1376 -190 1396 -135

rect 1502 -190 1525 -135

rect 1629 -190 1651 -135

rect 1758 -190 1778 -135

rect 1886 -190 1906 -135

rect 2012 -190 2035 -135

rect -58 -195 2122 -190

rect -58 -197 66 -195

rect -58 -217 -31 -197

rect -11 -217 6 -197

rect 26 -215 66 -197

rect 86 -197 134 -195

rect 86 -215 99 -197

rect 26 -217 99 -215

rect 119 -215 134 -197

rect 154 -215 186 -195

rect 206 -215 224 -195

rect 244 -197 579 -195

rect 244 -198 314 -197

rect 244 -215 268 -198

rect 119 -217 268 -215

rect -58 -218 268 -217

rect 288 -217 314 -198

rect 334 -198 395 -197

rect 334 -217 353 -198

rect 288 -218 353 -217

rect 373 -217 395 -198

rect 415 -217 442 -197

rect 462 -217 479 -197

rect 499 -217 527 -197

rect 547 -215 579 -197

rect 596 -197 644 -195

rect 596 -215 609 -197

rect 547 -217 609 -215

rect 629 -215 644 -197

rect 664 -215 696 -195

rect 716 -215 734 -195

rect 754 -197 1217 -195

rect 754 -198 824 -197

rect 754 -215 778 -198

rect 629 -217 778 -215

rect 373 -218 778 -217

rect 798 -217 824 -198

rect 844 -198 905 -197

rect 844 -217 863 -198

rect 798 -218 863 -217

rect 883 -217 905 -198

rect 925 -217 952 -197

rect 972 -217 989 -197

rect 1009 -217 1037 -197

rect 1057 -217 1120 -197

rect 1140 -217 1157 -197

rect 1177 -215 1217 -197

rect 1237 -197 1285 -195

rect 1237 -215 1250 -197

rect 1177 -217 1250 -215

rect 1270 -215 1285 -197

rect 1305 -215 1337 -195

rect 1357 -215 1375 -195

rect 1395 -197 1730 -195

rect 1395 -198 1465 -197

rect 1395 -215 1419 -198

rect 1270 -217 1419 -215

rect 883 -218 1419 -217

rect 1439 -217 1465 -198

rect 1485 -198 1546 -197

rect 1485 -217 1504 -198

rect 1439 -218 1504 -217

rect 1524 -217 1546 -198

rect 1566 -217 1593 -197

rect 1613 -217 1630 -197

rect 1650 -217 1678 -197

rect 1698 -215 1730 -197

rect 1747 -197 1795 -195

rect 1747 -215 1760 -197

rect 1698 -217 1760 -215

rect 1780 -215 1795 -197

rect 1815 -215 1847 -195

rect 1867 -215 1885 -195

rect 1905 -196 2122 -195

rect 1905 -197 2088 -196

rect 1905 -198 1975 -197

rect 1905 -215 1929 -198

rect 1780 -217 1929 -215

rect 1524 -218 1929 -217

rect 1949 -217 1975 -198

rect 1995 -198 2051 -197

rect 1995 -217 2014 -198

rect 1949 -218 2014 -217

rect 2034 -217 2051 -198

rect 2071 -216 2088 -197

rect 2108 -216 2122 -196

rect 2071 -217 2122 -216

rect 2034 -218 2122 -217

rect -58 -221 2122 -218

<< viali >>

rect -30 116 -10 136

rect 98 118 118 138

rect 221 117 241 137

rect 350 116 370 136

rect 481 116 501 136

rect 608 118 628 138

rect 731 117 751 137

rect 860 116 880 136

rect 991 116 1011 136

rect 1121 116 1141 136

rect 1249 118 1269 138

rect 1372 117 1392 137

rect 1501 116 1521 136

rect 1632 116 1652 136

rect 1759 118 1779 138

rect 1882 117 1902 137

rect 2011 116 2031 136

rect -26 -53 -6 -33

rect 2093 -50 2113 -30

rect -31 -217 -11 -197

rect 99 -217 119 -197

rect 224 -215 244 -195

rect 353 -218 373 -198

rect 479 -217 499 -197

rect 609 -217 629 -197

rect 734 -215 754 -195

rect 863 -218 883 -198

rect 989 -217 1009 -197

rect 1120 -217 1140 -197

rect 1250 -217 1270 -197

rect 1375 -215 1395 -195

rect 1504 -218 1524 -198

rect 1630 -217 1650 -197

rect 1760 -217 1780 -197

rect 1885 -215 1905 -195

rect 2014 -218 2034 -198

<< metal1 >>

rect -60 138 2123 142

rect -60 136 98 138

rect -60 116 -30 136

rect -10 118 98 136

rect 118 137 608 138

rect 118 118 221 137

rect -10 117 221 118

rect 241 136 608 137

rect 241 117 350 136

rect -10 116 350 117

rect 370 116 481 136

rect 501 118 608 136

rect 628 137 1249 138

rect 628 118 731 137

rect 501 117 731 118

rect 751 136 1249 137

rect 751 117 860 136

rect 501 116 860 117

rect 880 116 991 136

rect 1011 116 1121 136

rect 1141 118 1249 136

rect 1269 137 1759 138

rect 1269 118 1372 137

rect 1141 117 1372 118

rect 1392 136 1759 137

rect 1392 117 1501 136

rect 1141 116 1501 117

rect 1521 116 1632 136

rect 1652 118 1759 136

rect 1779 137 2123 138

rect 1779 118 1882 137

rect 1652 117 1882 118

rect 1902 136 2123 137

rect 1902 117 2011 136

rect 1652 116 2011 117

rect 2031 116 2123 136

rect -60 111 2123 116

rect -32 -32 2 -28

rect 2084 -30 2120 -26

rect 2084 -32 2093 -30

rect -32 -33 2093 -32

rect -32 -53 -26 -33

rect -6 -50 2093 -33

rect 2113 -50 2120 -30

rect -6 -52 2120 -50

rect -6 -53 2 -52

rect -32 -59 2 -53

rect 2084 -57 2120 -52

rect 1500 -190 1538 -189

rect -58 -195 2122 -190

rect -58 -197 224 -195

rect -58 -217 -31 -197

rect -11 -217 99 -197

rect 119 -215 224 -197

rect 244 -197 734 -195

rect 244 -198 479 -197

rect 244 -215 353 -198

rect 119 -217 353 -215

rect -58 -218 353 -217

rect 373 -217 479 -198

rect 499 -217 609 -197

rect 629 -215 734 -197

rect 754 -197 1375 -195

rect 754 -198 989 -197

rect 754 -215 863 -198

rect 629 -217 863 -215

rect 373 -218 863 -217

rect 883 -217 989 -198

rect 1009 -217 1120 -197

rect 1140 -217 1250 -197

rect 1270 -215 1375 -197

rect 1395 -197 1885 -195

rect 1395 -198 1630 -197

rect 1395 -215 1504 -198

rect 1270 -217 1504 -215

rect 883 -218 1504 -217

rect 1524 -217 1630 -198

rect 1650 -217 1760 -197

rect 1780 -215 1885 -197

rect 1905 -198 2122 -195

rect 1905 -215 2014 -198

rect 1780 -217 2014 -215

rect 1524 -218 2014 -217

rect 2034 -218 2122 -198

rect -58 -221 2122 -218

<< labels >>

flabel locali s -57 111 -20 140 0 FreeSans 80 0 0 0 VDD

port 0 nsew

flabel locali s -53 -219 -16 -190 0 FreeSans 80 0 0 0 GND

port 1 nsew

flabel locali s 2083 -56 2121 -27 0 FreeSans 80 0 0 0 OUT

port 2 nsew

<< end >>
