* SPICE3 file created from priority_encoder.ext - technology: sky130A
.include pshort.lib
.include nshort.lib
.option scale=0.01u

//.subckt priority_encoder VDD GND I0 I1 I2 I3 O0 O1
M1000 a_246_127# I1 a_246_n127# GND nshort_model.0 ad=4080 pd=262 as=2160 ps=134 w=80 l=18
M1001 a_976_n127# I3 GND GND nshort_model.0 ad=2160 pd=134 as=4080 ps=262 w=80 l=18
M1002 O0 a_610_n127# VDD VDD pshort_model.0 ad=4000 pd=258 as=4000 ps=258 w=77 l=18
M1003 a_464_n127# a_246_127# GND GND nshort_model.0 ad=4000 pd=260 as=4000 ps=260 w=80 l=18
M1004 VDD I1 a_246_127# VDD pshort_model.0 ad=3720 pd=250 as=2050 ps=130 w=76 l=18
M1005 a_610_n127# a_464_n127# GND GND nshort_model.0 ad=2160 pd=134 as=4080 ps=262 w=80 l=18
M1006 a_246_127# a_78_n127# VDD VDD pshort_model.0 ad=2050 pd=130 as=3720 ps=250 w=76 l=18
M1007 a_976_n127# I2 a_976_127# VDD pshort_model.0 ad=3720 pd=250 as=2050 ps=130 w=76 l=18
M1008 a_n71_n128# I0 GND GND nshort_model.0 ad=4000 pd=260 as=4000 ps=260 w=80 l=18
M1009 GND I2 a_976_n127# GND nshort_model.0 ad=4080 pd=262 as=2160 ps=134 w=80 l=18
M1010 a_610_n127# I3 a_610_127# VDD pshort_model.0 ad=3720 pd=250 as=2050 ps=130 w=76 l=18
M1011 O1 a_976_n127# GND GND nshort_model.0 ad=4000 pd=260 as=4000 ps=260 w=80 l=18
M1012 GND I3 a_610_n127# GND nshort_model.0 ad=4080 pd=262 as=2160 ps=134 w=80 l=18
M1013 a_976_127# I3 VDD VDD pshort_model.0 ad=2050 pd=130 as=3720 ps=250 w=76 l=18
M1014 O0 a_610_n127# GND GND nshort_model.0 ad=4000 pd=260 as=4000 ps=260 w=80 l=18
M1015 a_78_n127# I2 VDD VDD pshort_model.0 ad=4000 pd=258 as=4000 ps=258 w=77 l=18
M1016 a_464_n127# a_246_127# VDD VDD pshort_model.0 ad=4000 pd=258 as=4000 ps=258 w=77 l=18
M1017 a_610_127# a_464_n127# VDD VDD pshort_model.0 ad=2050 pd=130 as=3720 ps=250 w=76 l=18
M1018 a_78_n127# I2 GND GND nshort_model.0 ad=4000 pd=260 as=4000 ps=260 w=80 l=18
M1019 a_246_n127# a_78_n127# GND GND nshort_model.0 ad=2160 pd=134 as=4080 ps=262 w=80 l=18
M1020 a_n71_n128# I0 VDD VDD pshort_model.0 ad=4000 pd=258 as=4000 ps=258 w=77 l=18
M1021 O1 a_976_n127# VDD VDD pshort_model.0 ad=4000 pd=258 as=4000 ps=258 w=77 l=18

VDD VDD 0 5V
VSS VSS 0 0V
Va I0 0 5V
Vb I1 0 5V
Vc I2 0 5V
Vd I3 0 0V


C0 VDD I2 0.0586f
C1 a_78_n127# I2 0.18f
C2 a_610_n127# I2 0.0551f
C3 a_246_127# I2 0.0667f
C4 a_464_n127# VDD 0.359f
C5 a_464_n127# a_610_n127# 0.122f
C6 O1 VDD 0.165f
C7 VDD I0 0.0255f
C8 a_464_n127# a_246_127# 0.194f
C9 a_78_n127# I0 2.49e-20
C10 I2 a_610_127# 0.00282f
C11 O0 VDD 0.251f
C12 I2 a_976_127# 0.00282f
C13 a_610_n127# O0 0.126f
C14 a_78_n127# VDD 0.33f
C15 I2 a_246_n127# 0.00524f
C16 a_976_n127# I2 0.227f
C17 a_610_n127# VDD 0.314f
C18 a_246_127# VDD 0.453f
C19 a_78_n127# a_246_127# 0.0705f
C20 I2 I1 0.0134f
C21 I2 I3 0.493f
C22 O1 a_976_n127# 0.13f
C23 VDD a_610_127# 0.0218f
C24 a_610_n127# a_610_127# 0.0156f
C25 a_464_n127# I1 2.41e-19
C26 O0 a_976_n127# 0.0285f
C27 VDD a_976_127# 0.0218f
C28 a_464_n127# I3 0.0987f
C29 VDD a_976_n127# 0.307f
C30 I2 a_n71_n128# 0.0245f
C31 a_246_127# a_246_n127# 0.0129f
C32 O0 I3 0.0725f
C33 VDD I1 0.0242f
C34 VDD I3 0.14f
C35 a_78_n127# I1 0.0981f
C36 a_610_n127# I3 0.295f
C37 a_246_127# I1 0.102f
C38 I0 a_n71_n128# 0.0413f
C39 a_976_n127# a_976_127# 0.0159f
C40 a_464_n127# I2 0.0623f
C41 VDD a_n71_n128# 0.256f
C42 a_78_n127# a_n71_n128# 0.0361f
C43 O1 I2 0.0111f
C44 I2 I0 0.0419f
C45 a_976_n127# I3 0.0994f
C46 O0 I2 0.0382f
C47 O1 GND 0.42f
C48 O0 GND 0.384f
C49 I3 GND 0.834f
C50 I1 GND 0.283f
C51 I2 GND 1.65f
C52 I0 GND 0.348f
C53 VDD GND 6.16f
C54 a_246_n127# GND 0.0226f 
C55 a_n71_n128# GND 0.426f 
C56 a_976_n127# GND 0.858f 
C57 a_610_n127# GND 0.821f 
C58 a_464_n127# GND 0.766f
C59 a_246_127# GND 0.766f 
C60 a_78_n127# GND 0.788f 
.ends
.tran 1n 100n
.control
run
.endc
.end
