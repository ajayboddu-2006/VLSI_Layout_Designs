magic
tech sky130A
timestamp 1736957124
<< nwell >>
rect -88 52 88 199
<< nmos >>
rect -2 -38 13 13
<< pmos >>
rect -2 71 13 121
<< ndiff >>
rect -41 5 -2 13
rect -41 -30 -34 5
rect -16 -30 -2 5
rect -41 -38 -2 -30
rect 13 6 55 13
rect 13 -32 27 6
rect 45 -32 55 6
rect 13 -38 55 -32
<< pdiff >>
rect -39 114 -2 121
rect -39 79 -32 114
rect -14 79 -2 114
rect -39 71 -2 79
rect 13 114 55 121
rect 13 76 27 114
rect 47 76 55 114
rect 13 71 55 76
<< ndiffc >>
rect -34 -30 -16 5
rect 27 -32 45 6
<< pdiffc >>
rect -32 79 -14 114
rect 27 76 47 114
<< psubdiff >>
rect -80 -69 95 -66
rect -80 -70 66 -69
rect -80 -87 -2 -70
rect 15 -87 32 -70
rect 49 -86 66 -70
rect 83 -86 95 -69
rect 49 -87 95 -86
rect -80 -91 95 -87
<< nsubdiff >>
rect -67 178 62 181
rect -67 161 -3 178
rect 15 161 32 178
rect 50 161 62 178
rect -67 156 62 161
<< psubdiffcont >>
rect -2 -87 15 -70
rect 32 -87 49 -70
rect 66 -86 83 -69
<< nsubdiffcont >>
rect -3 161 15 178
rect 32 161 50 178
<< poly >>
rect -2 121 13 140
rect -2 49 13 71
rect -23 34 13 49
rect -2 13 13 34
rect -2 -51 13 -38
<< locali >>
rect -89 178 86 181
rect -89 161 -77 178
rect -60 161 -34 178
rect -17 161 -3 178
rect 15 161 32 178
rect 50 161 86 178
rect -89 156 86 161
rect -35 121 -12 156
rect -39 114 -8 121
rect -39 79 -32 114
rect -14 79 -8 114
rect -39 71 -8 79
rect 19 114 55 121
rect 19 76 27 114
rect 47 76 55 114
rect 19 71 55 76
rect 25 50 49 71
rect 25 30 60 50
rect 25 13 49 30
rect -41 5 -8 13
rect -41 -30 -34 5
rect -16 -30 -8 5
rect -41 -38 -8 -30
rect 19 6 55 13
rect 19 -32 27 6
rect 45 -32 55 6
rect 19 -38 55 -32
rect -36 -66 -13 -38
rect -80 -69 95 -66
rect -80 -70 66 -69
rect -80 -87 -72 -70
rect -55 -87 -34 -70
rect -17 -87 -2 -70
rect 15 -87 32 -70
rect 49 -86 66 -70
rect 83 -86 95 -69
rect 49 -87 95 -86
rect -80 -91 95 -87
<< viali >>
rect -77 161 -60 178
rect -34 161 -17 178
rect -72 -87 -55 -70
rect -34 -87 -17 -70
<< metal1 >>
rect -89 178 86 181
rect -89 161 -77 178
rect -60 161 -34 178
rect -17 161 86 178
rect -89 156 86 161
rect -80 -70 95 -66
rect -80 -87 -72 -70
rect -55 -87 -34 -70
rect -17 -87 95 -70
rect -80 -91 95 -87
<< labels >>
flabel metal1 s -87 159 -66 177 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel metal1 s -76 -87 -55 -69 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel poly s -24 34 -3 52 0 FreeSans 80 0 0 0 IN
port 2 nsew
flabel locali s 27 31 48 49 0 FreeSans 80 0 0 0 OUT
port 3 nsew
<< end >>
