magic

tech sky130A

timestamp 1737028004

<< nwell >>

rect -86 148 281 290

rect 114 141 281 148

<< nmos >>

rect -27 34 -12 82

rect 24 34 39 82

rect 212 35 227 80

<< pmos >>

rect -27 166 -12 211

rect 24 166 39 211

rect 212 164 227 212

<< ndiff >>

rect -64 74 -27 82

rect -64 42 -55 74

rect -34 42 -27 74

rect -64 34 -27 42

rect -12 34 24 82

rect 39 74 78 82

rect 39 42 49 74

rect 70 42 78 74

rect 39 34 78 42

rect 182 72 212 80

rect 182 43 189 72

rect 206 43 212 72

rect 182 35 212 43

rect 227 72 257 80

rect 227 43 236 72

rect 253 43 257 72

rect 227 35 257 43

<< pdiff >>

rect -62 204 -27 211

rect -62 173 -54 204

rect -37 173 -27 204

rect -62 166 -27 173

rect -12 204 24 211

rect -12 173 -2 204

rect 15 173 24 204

rect -12 166 24 173

rect 39 204 72 211

rect 39 173 48 204

rect 65 173 72 204

rect 39 166 72 173

rect 185 204 212 212

rect 185 172 189 204

rect 206 172 212 204

rect 185 164 212 172

rect 227 204 255 212

rect 227 172 234 204

rect 251 172 255 204

rect 227 164 255 172

<< ndiffc >>

rect -55 42 -34 74

rect 49 42 70 74

rect 189 43 206 72

rect 236 43 253 72

<< pdiffc >>

rect -54 173 -37 204

rect -2 173 15 204

rect 48 173 65 204

rect 189 172 206 204

rect 234 172 251 204

<< psubdiff >>

rect -94 -5 285 -2

rect -94 -22 -80 -5

rect -63 -6 78 -5

rect -63 -22 -25 -6

rect -94 -23 -25 -22

rect -8 -23 9 -6

rect 26 -23 44 -6

rect 61 -22 78 -6

rect 95 -6 255 -5

rect 95 -22 112 -6

rect 61 -23 112 -22

rect 129 -23 146 -6

rect 163 -23 218 -6

rect 235 -22 255 -6

rect 272 -22 285 -5

rect 235 -23 285 -22

rect -94 -27 285 -23

<< nsubdiff >>

rect -68 269 260 272

rect -68 268 36 269

rect -68 251 -34 268

rect -17 251 0 268

rect 17 252 36 268

rect 53 252 83 269

rect 100 252 117 269

rect 134 252 152 269

rect 169 252 231 269

rect 248 252 260 269

rect 17 251 260 252

rect -68 247 260 251

<< psubdiffcont >>

rect -80 -22 -63 -5

rect -25 -23 -8 -6

rect 9 -23 26 -6

rect 44 -23 61 -6

rect 78 -22 95 -5

rect 112 -23 129 -6

rect 146 -23 163 -6

rect 218 -23 235 -6

rect 255 -22 272 -5

<< nsubdiffcont >>

rect -34 251 -17 268

rect 0 251 17 268

rect 36 252 53 269

rect 83 252 100 269

rect 117 252 134 269

rect 152 252 169 269

rect 231 252 248 269

<< poly >>

rect -27 211 -12 233

rect 24 211 39 233

rect 212 212 227 230

rect -89 137 -58 145

rect -89 120 -80 137

rect -63 135 -58 137

rect -27 135 -12 166

rect -63 120 -12 135

rect -89 112 -58 120

rect -27 82 -12 120

rect 24 143 39 166

rect 75 143 114 149

rect 24 141 114 143

rect 24 124 87 141

rect 104 124 114 141

rect 24 82 39 124

rect 75 117 114 124

rect 152 122 185 127

rect 212 122 227 164

rect 152 120 227 122

rect 152 103 160 120

rect 177 103 227 120

rect 152 97 185 103

rect 212 80 227 103

rect -27 14 -12 34

rect 24 14 39 34

rect 212 13 227 35

<< polycont >>

rect -80 120 -63 137

rect 87 124 104 141

rect 160 103 177 120

<< locali >>

rect -86 269 280 272

rect -86 252 -63 269

rect -46 268 36 269

rect -46 252 -34 268

rect -86 251 -34 252

rect -17 251 0 268

rect 17 252 36 268

rect 53 252 55 269

rect 72 252 83 269

rect 100 252 117 269

rect 134 252 152 269

rect 169 252 185 269

rect 202 252 231 269

rect 248 252 280 269

rect 17 251 280 252

rect -86 247 280 251

rect -62 211 -45 247

rect 55 211 72 247

rect 185 212 202 247

rect -62 204 -29 211

rect -62 173 -54 204

rect -37 173 -29 204

rect -62 166 -29 173

rect -10 204 23 211

rect -10 173 -2 204

rect 15 173 23 204

rect -10 166 23 173

rect 40 204 73 211

rect 40 173 48 204

rect 65 173 73 204

rect 40 166 73 173

rect 185 204 210 212

rect 185 172 189 204

rect 206 172 210 204

rect -89 137 -58 145

rect -97 120 -80 137

rect -63 120 -58 137

rect -2 131 15 166

rect 185 164 210 172

rect 229 204 255 212

rect 229 172 234 204

rect 251 172 255 204

rect 229 164 255 172

rect 75 141 114 149

rect -89 112 -58 120

rect -15 124 24 131

rect -15 107 -5 124

rect 13 116 24 124

rect 75 124 87 141

rect 104 124 120 141

rect 235 130 254 164

rect 75 121 120 124

rect 75 117 114 121

rect 152 120 185 127

rect 13 107 58 116

rect -15 99 58 107

rect 41 82 58 99

rect 152 103 160 120

rect 177 103 185 120

rect 152 97 185 103

rect 235 111 268 130

rect -64 74 -28 82

rect -64 42 -55 74

rect -34 42 -28 74

rect -64 34 -28 42

rect 41 74 78 82

rect 235 80 254 111

rect 41 42 49 74

rect 70 42 78 74

rect 41 34 78 42

rect 182 72 211 80

rect 182 43 189 72

rect 206 43 211 72

rect 182 35 211 43

rect 228 72 257 80

rect 228 43 236 72

rect 253 43 257 72

rect 228 35 257 43

rect -57 -2 -39 34

rect 186 -2 204 35

rect -94 -5 285 -2

rect -94 -22 -80 -5

rect -63 -6 78 -5

rect -63 -22 -56 -6

rect -94 -23 -56 -22

rect -39 -23 -25 -6

rect -8 -23 9 -6

rect 26 -23 44 -6

rect 61 -22 78 -6

rect 95 -6 255 -5

rect 95 -22 112 -6

rect 61 -23 112 -22

rect 129 -23 146 -6

rect 163 -23 185 -6

rect 202 -23 218 -6

rect 235 -22 255 -6

rect 272 -22 285 -5

rect 235 -23 285 -22

rect -94 -27 285 -23

<< viali >>

rect -63 252 -46 269

rect 55 252 72 269

rect 185 252 202 269

rect -5 107 13 124

rect 160 103 177 120

rect -56 -23 -39 -6

rect 185 -23 202 -6

<< metal1 >>

rect -86 269 280 272

rect -86 252 -63 269

rect -46 252 55 269

rect 72 252 185 269

rect 202 252 280 269

rect -86 247 280 252

rect -15 124 24 131

rect -15 107 -5 124

rect 13 116 24 124

rect 152 120 185 128

rect 152 116 160 120

rect 13 107 160 116

rect -15 103 160 107

rect 177 103 185 120

rect -15 99 185 103

rect 152 97 185 99

rect -94 -6 285 -2

rect -94 -23 -56 -6

rect -39 -23 185 -6

rect 202 -23 285 -6

rect -94 -27 285 -23

<< labels >>

flabel space -89 248 -62 269 0 FreeSans 80 0 0 0 VDD

port 0 nsew

flabel locali -88 115 -61 136 0 FreeSans 80 0 0 0 IN1

port 2 nsew

flabel metal1 -93 -25 -66 -4 0 FreeSans 80 0 0 0 GND

port 1 nsew

flabel locali 81 123 108 144 0 FreeSans 80 0 0 0 IN2

port 3 nsew

flabel locali s 237 112 264 133 0 FreeSans 80 0 0 0 OUT

port 4 nsew

<< end >>
