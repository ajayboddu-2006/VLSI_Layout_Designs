* SPICE3 file created from Full_Adder.ext - technology: sky130A
.include pshort.lib
.include nshort.lib
.option scale=0.01u

//.subckt Full_Adder VDD GND A B Cin SUM COUT
M1000 a_654_n141# a_494_9# VDD VDD pshort_model.0 ad=1620 pd=162 as=1490 ps=156 w=45 l=15
M1001 a_494_9# B a_494_n141# GND nshort_model.0 ad=1540 pd=158 as=770 ps=79u w=44 l=15
M1002 a_1654_n141# a_654_n141# GND GND nshort_model.0 ad=814 pd=81u as=1500 ps=156 w=44 l=15
M1003 a_n117_n141# A VDD VDD pshort_model.0 ad=1670 pd=164 as=1620 ps=162 w=45 l=15
M1004 a_1380_9# a_382_n141# VDD VDD pshort_model.0 ad=787 pd=80u as=1580 ps=160 w=45 l=15
M1005 a_n3_n147# B VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1006 a_949_9# a_382_n141# a_1049_n146# VDD pshort_model.0 ad=1670 pd=164 as=770 ps=79u w=44 l=15
M1007 COUT a_1654_n141# VDD VDD pshort_model.0 ad=1670 pd=164 as=1620 ps=162 w=45 l=15
M1008 GND A a_213_n146# GND nshort_model.0 ad=1410 pd=152 as=770 ps=79u w=44 l=15
M1009 a_1380_9# Cin a_1380_n141# GND nshort_model.0 ad=1540 pd=158 as=770 ps=79u w=44 l=15
M1010 COUT a_1654_n141# GND GND nshort_model.0 ad=1510 pd=156 as=1510 ps=156 w=42 l=15
M1011 a_163_n146# a_n3_n147# a_63_9# VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1012 GND a_382_n141# a_1099_n146# GND nshort_model.0 ad=1410 pd=152 as=770 ps=79u w=44 l=15
M1013 a_999_n146# a_769_n141# GND GND nshort_model.0 ad=770 pd=79u as=1500 ps=156 w=44 l=15
M1014 GND a_1540_n141# a_1654_n141# GND nshort_model.0 ad=1500 pd=156 as=814 ps=81u w=44 l=15
M1015 a_63_9# B VDD VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1016 a_163_n146# B a_113_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1017 VDD Cin a_1380_9# VDD pshort_model.0 ad=1580 pd=160 as=787 ps=80u w=45 l=15
M1018 a_883_n147# Cin GND GND nshort_model.0 ad=1580 pd=160 as=1580 ps=160 w=45 l=15
M1019 VDD a_n117_n141# a_63_9# VDD pshort_model.0 ad=770 pd=79u as=1540 ps=158 w=44 l=15
M1020 a_1654_9# a_654_n141# VDD VDD pshort_model.0 ad=832 pd=82u as=1620 ps=162 w=45 l=15
M1021 a_1049_n146# Cin a_999_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1022 a_494_9# A VDD VDD pshort_model.0 ad=787 pd=80u as=1580 ps=160 w=45 l=15
M1023 a_654_n141# a_494_9# GND GND nshort_model.0 ad=1500 pd=156 as=1450 ps=154 w=44 l=15
M1024 SUM a_1049_n146# VDD VDD pshort_model.0 ad=1580 pd=160 as=1530 ps=158 w=45 l=15
M1025 a_63_9# A a_163_n146# VDD pshort_model.0 ad=1670 pd=164 as=770 ps=79u w=44 l=15
M1026 a_883_n147# Cin VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1027 a_1540_n141# a_1380_9# VDD VDD pshort_model.0 ad=1620 pd=162 as=1490 ps=156 w=45 l=15
M1028 a_1540_n141# a_1380_9# GND GND nshort_model.0 ad=1500 pd=156 as=1450 ps=154 w=44 l=15
M1029 a_769_n141# a_382_n141# VDD VDD pshort_model.0 ad=1670 pd=164 as=1620 ps=162 w=45 l=15
M1030 a_n117_n141# A GND GND nshort_model.0 ad=1510 pd=156 as=1510 ps=156 w=42 l=15
M1031 a_1654_n141# a_1540_n141# a_1654_9# VDD pshort_model.0 ad=1620 pd=162 as=832 ps=82u w=45 l=15
M1032 a_1049_n146# a_883_n147# a_949_9# VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1033 a_113_n146# a_n117_n141# GND GND nshort_model.0 ad=770 pd=79u as=1500 ps=156 w=44 l=15
M1034 a_494_n141# A GND GND nshort_model.0 ad=770 pd=79u as=1450 ps=154 w=44 l=15
M1035 a_n3_n147# B GND GND nshort_model.0 ad=1580 pd=160 as=1580 ps=160 w=45 l=15
M1036 VDD B a_494_9# VDD pshort_model.0 ad=1580 pd=160 as=787 ps=80u w=45 l=15
M1037 a_382_n141# a_163_n146# GND GND nshort_model.0 ad=1500 pd=156 as=1500 ps=156 w=44 l=15
M1038 a_213_n146# a_n3_n147# a_163_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1039 a_1380_n141# a_382_n141# GND GND nshort_model.0 ad=770 pd=79u as=1450 ps=154 w=44 l=15
M1040 VDD a_769_n141# a_949_9# VDD pshort_model.0 ad=770 pd=79u as=1540 ps=158 w=44 l=15
M1041 a_949_9# Cin VDD VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1042 a_769_n141# a_382_n141# GND GND nshort_model.0 ad=1510 pd=156 as=1510 ps=156 w=42 l=15
M1043 SUM a_1049_n146# GND GND nshort_model.0 ad=1500 pd=156 as=1500 ps=156 w=44 l=15
M1044 a_382_n141# a_163_n146# VDD VDD pshort_model.0 ad=1580 pd=160 as=1530 ps=158 w=45 l=15
M1045 a_1099_n146# a_883_n147# a_1049_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15

VDD VDD 0 5V
VSS VSS 0 0V
Va A VSS PULSE(0 5V 0 0.1ns 0.1ns 8ns 16ns)
Vb B VSS PULSE(0 5V 0 0.1ns 0.1ns 15ns 30ns)
Vc Cin VSS PULSE(0 5V 0 0.1ns 0.1ns 7ns 14ns)

C0 a_654_n141# A 7.96e-19
C1 a_654_n141# VDD 0.257f
C2 a_163_n146# a_213_n146# 0.00731f
C3 a_382_n141# B 0.00947f
C4 a_382_n141# a_1049_n146# 0.251f
C5 VDD a_494_n141# 5.82e-21
C6 a_769_n141# a_494_9# 9.99e-20
C7 a_163_n146# a_63_9# 0.228f
C8 a_1654_n141# COUT 0.107f
C9 a_382_n141# a_654_n141# 0.319f
C10 a_163_n146# a_113_n146# 0.00374f
C11 a_1380_9# VDD 0.264f
C12 a_769_n141# a_949_9# 0.0121f
C13 a_382_n141# a_494_n141# 0.00172f
C14 a_494_9# A 0.0187f
C15 a_1540_n141# a_654_n141# 0.26f
C16 a_1049_n146# a_883_n147# 0.171f
C17 a_494_9# VDD 0.26f
C18 a_382_n141# a_1380_9# 0.0706f
C19 a_654_n141# a_883_n147# 0.0165f
C20 VDD a_1380_n141# 1.69e-19
C21 a_769_n141# Cin 0.155f
C22 a_n117_n141# a_n3_n147# 0.229f
C23 a_1654_n141# VDD 0.145f
C24 a_1654_n141# a_1654_9# 0.00403f
C25 a_949_9# VDD 0.551f
C26 a_1540_n141# a_1380_9# 0.0655f
C27 a_382_n141# a_494_9# 0.13f
C28 a_63_9# A 0.0136f
C29 a_63_9# VDD 0.551f
C30 a_382_n141# a_949_9# 0.423f
C31 a_n117_n141# B 0.158f
C32 VDD Cin 0.0466f
C33 a_1049_n146# SUM 0.077f
C34 a_1049_n146# a_999_n146# 0.00374f
C35 a_382_n141# a_63_9# 0.00219f
C36 a_654_n141# SUM 0.0115f
C37 a_1654_n141# a_1540_n141# 0.202f
C38 a_654_n141# a_999_n146# 0.00132f
C39 a_382_n141# Cin 0.141f
C40 a_949_9# a_883_n147# 0.149f
C41 a_163_n146# A 0.105f
C42 a_1380_9# SUM 0.0265f
C43 a_1540_n141# Cin 7.94e-19
C44 a_163_n146# VDD 0.0681f
C45 a_883_n147# Cin 0.152f
C46 a_n3_n147# B 0.152f
C47 COUT VDD 0.115f
C48 a_382_n141# a_163_n146# 0.0608f
C49 a_769_n141# VDD 0.198f
C50 a_382_n141# a_1099_n146# 0.0017f
C51 a_949_9# SUM 0.00219f
C52 a_n117_n141# a_63_9# 0.0253f
C53 a_382_n141# a_769_n141# 0.355f
C54 VDD A 0.042f
C55 a_1540_n141# COUT 1.85e-19
C56 a_654_n141# B 0.00144f
C57 a_1049_n146# a_654_n141# 0.0263f
C58 SUM Cin 2.46e-19
C59 VDD a_1654_9# 0.00956f
C60 a_382_n141# A 0.0169f
C61 a_769_n141# a_883_n147# 0.22f
C62 a_382_n141# VDD 0.71f
C63 a_654_n141# a_1380_9# 0.0671f
C64 a_n117_n141# a_163_n146# 0.0157f
C65 a_1540_n141# VDD 0.294f
C66 a_1540_n141# a_1654_9# 0.00395f
C67 a_494_9# B 0.0812f
C68 a_63_9# a_n3_n147# 0.163f
C69 a_n3_n147# a_113_n146# 0.00282f
C70 a_883_n147# VDD 0.186f
C71 a_654_n141# a_494_9# 0.0782f
C72 a_382_n141# a_1540_n141# 2.11e-19
C73 a_1049_n146# a_949_9# 0.211f
C74 a_654_n141# a_1380_n141# 0.00133f
C75 a_494_9# a_494_n141# 0.00699f
C76 a_1654_n141# a_654_n141# 0.056f
C77 a_63_9# B 0.0137f
C78 a_382_n141# a_883_n147# 0.17f
C79 a_654_n141# a_949_9# 0.0129f
C80 a_1049_n146# Cin 0.0107f
C81 a_1380_9# a_1380_n141# 0.00699f
C82 a_n117_n141# A 0.025f
C83 a_163_n146# a_n3_n147# 0.171f
C84 a_654_n141# Cin 0.0123f
C85 a_949_9# a_1380_9# 1.36e-19
C86 a_n117_n141# VDD 0.238f
C87 SUM VDD 0.178f
C88 a_1380_9# Cin 0.0812f
C89 a_382_n141# SUM 0.083f
C90 a_382_n141# a_999_n146# 0.0017f
C91 a_163_n146# B 0.0107f
C92 a_494_9# a_63_9# 1.36e-19
C93 a_1049_n146# a_1099_n146# 0.00731f
C94 a_654_n141# a_1099_n146# 0.00132f
C95 a_n3_n147# A 0.096f
C96 a_1049_n146# a_769_n141# 0.0157f
C97 a_63_9# a_213_n146# 0.00134f
C98 a_654_n141# COUT 1.16e-19
C99 a_883_n147# SUM 1.16e-19
C100 a_883_n147# a_999_n146# 0.00282f
C101 a_n3_n147# VDD 0.188f
C102 a_949_9# Cin 0.0111f
C103 a_769_n141# a_654_n141# 0.116f
C104 a_63_9# a_113_n146# 0.00134f
C105 a_382_n141# a_n3_n147# 4.98e-19
C106 A B 0.127f
C107 VDD B 0.0463f
C108 a_1049_n146# VDD 0.0721f
C109 COUT GND 0.254f
C110 SUM GND 0.237f
C111 Cin GND 0.511f
C112 B GND 0.511f
C113 A GND 0.578f
C114 VDD GND 7.18f
C115 a_1380_n141# GND 0.0088f **FLOATING
C116 a_1099_n146# GND 0.00892f **FLOATING
C117 a_999_n146# GND 0.00892f **FLOATING
C118 a_494_n141# GND 0.0088f **FLOATING
C119 a_213_n146# GND 0.00892f **FLOATING
C120 a_113_n146# GND 0.00892f **FLOATING
C121 a_1654_9# GND 1.22e-19 **FLOATING
C122 a_949_9# GND 0.0657f **FLOATING
C123 a_1654_n141# GND 0.704f **FLOATING
C124 a_1540_n141# GND 0.459f **FLOATING
C125 a_1380_9# GND 0.52f **FLOATING
C126 a_1049_n146# GND 0.561f **FLOATING
C127 a_883_n147# GND 0.479f **FLOATING
C128 a_769_n141# GND 0.687f **FLOATING
C129 a_654_n141# GND 1.38f **FLOATING
C130 a_63_9# GND 0.135f **FLOATING
C131 a_382_n141# GND 1.48f **FLOATING
C132 a_494_9# GND 0.525f **FLOATING
C133 a_163_n146# GND 0.578f **FLOATING
C134 a_n3_n147# GND 0.481f **FLOATING
C135 a_n117_n141# GND 0.746f **FLOATING
//.ends
.tran 1n 40n
.control
run
.endc
.end
