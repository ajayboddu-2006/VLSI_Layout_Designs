* SPICE3 file created from MUX_4X1.ext - technology: sky130A

.include pshort.lib
.include nshort.lib

.option scale=0.01u

//.subckt MUX_4X1 VDD GND I0 I1 I2 I3 S0 S1 OUT
M1000 a_373_267# S0 a_193_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1001 a_193_27# a_n240_27# a_133_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1002 a_15_27# I0 GND GND nmos_model.0 ad=1310 pd=104 as=2620 ps=208 w=61 l=15
M1003 a_253_27# S1 a_193_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1004 a_n113_27# S1 VDD VDD pmos_model.0 ad=2580 pd=206 as=2520 ps=204 w=60 l=15
M1005 VDD a_n113_27# a_15_267# VDD pmos_model.0 ad=1370 pd=106 as=1310 ps=104 w=61 l=15
M1006 a_193_267# I1 a_15_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1007 a_n240_27# S0 GND GND nmos_model.0 ad=2480 pd=202 as=2540 ps=204 w=59 l=15
M1008 GND I1 a_253_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1009 a_373_27# I2 GND GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1010 a_15_267# I0 VDD VDD pmos_model.0 ad=1310 pd=104 as=2620 ps=208 w=61 l=15
M1011 a_373_267# S1 a_133_27# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1012 a_73_27# a_n113_27# a_15_27# GND nmos_model.0 ad=1370 pd=106 as=1310 ps=104 w=61 l=15
M1013 a_433_27# a_n113_27# a_373_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1014 a_133_27# S0 a_433_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1015 a_553_27# S0 a_133_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1016 a_613_27# S1 a_553_27# GND nmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1017 GND I3 a_613_27# GND nmos_model.0 ad=2750 pd=212 as=1370 ps=106 w=61 l=15
M1018 a_15_267# a_n240_27# VDD VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1019 a_n240_27# S0 VDD VDD pmos_model.0 ad=2580 pd=206 as=2520 ps=204 w=60 l=15
M1020 a_193_267# a_n113_27# a_373_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1021 a_15_267# S1 a_193_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1022 a_n113_27# S1 GND GND nmos_model.0 ad=2540 pd=204 as=2540 ps=204 w=59 l=15
M1023 a_133_27# S0 a_373_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1024 OUT a_133_27# GND GND nmos_model.0 ad=2680 pd=210 as=2680 ps=210 w=61 l=15
M1025 a_373_267# I2 a_193_267# VDD pmos_model.0 ad=1370 pd=106 as=1370 ps=106 w=61 l=15
M1026 OUT a_133_27# VDD VDD pmos_model.0 ad=2750 pd=212 as=2750 ps=212 w=61 l=15
M1027 a_193_267# a_n240_27# a_15_267# VDD pmos_model.0 ad=1.37n pd=0.106m as=1.37n ps=0.106m w=61 l=15
M1028 a_133_27# I3 a_373_267# VDD pmos_model.0 ad=2.75n pd=0.212m as=1.37n ps=0.106m w=61 l=15
M1029 a_133_27# a_n240_27# a_73_27# GND nmos_model.0 ad=1.37n pd=0.106m as=1.37n ps=0.106m w=61 l=15

VDD VDD 0 5V
VSS VSS 0 0V
Va I0 PULSE(0 5V 0 0.1ns 0.1ns 2.5ns 5ns)
Va I1 PULSE(0 5V 0 0.1ns 0.1ns 5ns 10ns)
Va I2 PULSE(0 5V 0 0.1ns 0.1ns 10ns 20ns)
Va I3 PULSE(0 5V 0 0.1ns 0.1ns 20ns 40ns)
Va S0 PULSE(0 5V 0 0.1ns 0.1ns 50ns 100ns)
Va S1 PULSE(0 5V 0 0.1ns 0.1ns 25ns 50ns)

C0 a_15_27# a_133_27# 0.00445f
C1 a_133_27# a_373_267# 0.516f
C2 a_613_27# a_373_267# 7.9e-19
C3 a_133_27# a_n113_27# 0.0993f
C4 I1 a_15_267# 0.00797f
C5 I1 VDD 0.00349f
C6 a_253_27# a_n113_27# 0.00444f
C7 a_613_27# a_133_27# 0.00805f
C8 a_193_267# a_433_27# 6.61e-19
C9 S0 a_n240_27# 0.0391f
C10 I3 a_193_267# 1.47e-19
C11 S0 S1 0.182f
C12 I1 a_373_267# 0.00179f
C13 a_253_27# a_133_27# 0.00805f
C14 I1 a_n113_27# 0.019f
C15 a_n240_27# a_193_267# 0.0336f
C16 I2 a_193_267# 0.0225f
C17 OUT I3 1.53e-19
C18 a_193_267# S1 0.0225f
C19 I1 a_133_27# 0.0118f
C20 I3 S1 0.128f
C21 I2 a_n240_27# 3.09e-19
C22 a_n240_27# S1 0.166f
C23 VDD S0 0.0332f
C24 a_15_267# a_193_267# 0.511f
C25 a_373_27# a_n113_27# 0.0045f
C26 I0 a_n240_27# 0.0187f
C27 I0 S1 0.0511f
C28 VDD a_193_267# 0.256f
C29 a_n113_27# a_193_27# 0.00444f
C30 a_373_27# a_133_27# 0.00805f
C31 S0 a_373_267# 0.0327f
C32 S0 a_n113_27# 0.134f
C33 OUT VDD 0.142f
C34 a_133_27# a_193_27# 0.00994f
C35 a_193_267# a_373_267# 0.511f
C36 a_193_267# a_n113_27# 0.0674f
C37 I3 VDD 0.00869f
C38 S0 a_133_27# 0.076f
C39 a_n240_27# a_15_267# 0.153f
C40 I2 a_15_267# 0.00179f
C41 a_15_267# S1 0.0163f
C42 OUT a_373_267# 0.00112f
C43 I0 a_15_267# 0.00797f
C44 VDD a_n240_27# 0.451f
C45 I2 VDD 0.00347f
C46 a_193_267# a_133_27# 0.00303f
C47 VDD S1 0.0305f
C48 a_n113_27# a_433_27# 8.4e-19
C49 I3 a_373_267# 0.00797f
C50 I0 VDD 0.0182f
C51 OUT a_133_27# 0.092f
C52 a_133_27# a_433_27# 0.00994f
C53 I2 a_373_267# 0.00797f
C54 a_n240_27# a_n113_27# 0.591f
C55 I2 a_n113_27# 0.152f
C56 S1 a_373_267# 0.0163f
C57 a_n113_27# S1 0.0576f
C58 I3 a_133_27# 0.0915f
C59 I0 a_n113_27# 0.163f
C60 I1 a_193_267# 0.0224f
C61 a_n240_27# a_133_27# 0.0369f
C62 I2 a_133_27# 0.0122f
C63 a_133_27# S1 0.0585f
C64 VDD a_15_267# 0.583f
C65 I0 a_133_27# 0.00187f
C66 a_15_27# a_15_267# 5.93e-19
C67 a_15_267# a_373_267# 0.0358f
C68 a_15_267# a_n113_27# 0.0425f
C69 a_73_27# a_n113_27# 0.00448f
C70 I1 a_n240_27# 6.87e-19
C71 I1 I2 0.128f
C72 I1 S1 0.128f
C73 VDD a_373_267# 0.173f
C74 VDD a_n113_27# 0.219f
C75 a_553_27# a_133_27# 0.0147f
C76 a_15_267# a_133_27# 0.0466f
C77 a_73_27# a_133_27# 0.00651f
C78 VDD a_133_27# 0.117f
C79 a_15_27# a_n113_27# 0.00429f
C80 a_n113_27# a_373_267# 0.0344f
C81 S0 a_193_267# 0.0124f
C82 OUT GND 0.418f
C83 I3 GND 0.279f
C84 I2 GND 0.239f
C85 I1 GND 0.241f
C86 I0 GND 0.273f
C87 S1 GND 0.821f
C88 S0 GND 0.841f
C89 VDD GND 6.27f
C90 a_613_27# GND 0.0143f **FLOATING
C91 a_553_27# GND 0.0125f **FLOATING
C92 a_433_27# GND 0.0125f **FLOATING
C93 a_373_27# GND 0.0143f **FLOATING
C94 a_253_27# GND 0.0143f **FLOATING
C95 a_193_27# GND 0.0125f **FLOATING
C96 a_73_27# GND 0.0125f **FLOATING
C97 a_15_27# GND 0.0137f **FLOATING
C98 a_373_267# GND 0.133f **FLOATING
C99 a_193_267# GND 0.112f **FLOATING
C100 a_15_267# GND 0.124f **FLOATING
C101 a_133_27# GND 1.41f **FLOATING
C102 a_n240_27# GND 1.11f **FLOATING
C103 a_n113_27# GND 1.17f **FLOATING
//.ends
.tran 1n 100n
.control
run
.endc
.end 
