
* SPICE3 file created from AND.ext - technology: sky130A



.option scale=0.01u

.include pshort.lib

.include nshort.lib

//.subckt AND GND IN1 IN2 OUT



M1000 a_n12_166# IN1 w_n86_148# w_n86_148# pmos_model.0 ad=8100 pd=81u as=1580 ps=160 w=45 l=15

M1001 w_n86_148# IN2 a_n12_166# w_n86_148# pmos_model.0 ad=1490 pd= as=8100 ps=81u w=45 l=15

M1002 OUT a_n12_166# w_n86_148# w_n86_148# pmos_model.0 ad=1340 pd=152 as=1300 ps=150 w=48 l=15

M1003 a_n12_166# IN2 a_n12_34# GND nmos_model.0 ad=1870 pd=174 as=864 ps=84u w=48 l=15

M1004 a_n12_34# IN1 GND GND nmos_model.0 ad=864 pd=84u as=1780 ps=170 w=48 l=15

M1005 OUT a_n12_166# GND GND nmos_model.0 ad=1350 pd=150 as=1350 ps=150 w=45 l=15



VDD VDD 0 3.3V

VSS VSS 0 0V

Va IN1 VSS PULSE(0 3.3V 0 0.1ns  0.1ns 2ns 4ns)

Va IN2 VSS PULSE(0 3.3V 0 0.1ns  0.1ns 3ns 6ns)



C0 w_n86_148# IN2 0.0409f

C1 w_n86_148# a_n12_166# 0.335f

C2 w_n86_148# IN1 0.0382f

C3 w_n86_148# OUT 0.121f

C4 IN2 a_n12_166# 0.129f

C5 IN2 IN1 0.0805f

C6 IN1 a_n12_166# 0.0498f

C7 IN2 OUT 0.00623f

C8 OUT a_n12_166# 0.048f

C9 a_n12_166# a_n12_34# 0.0105f

C10 OUT GND 0.259f

C11 IN2 GND 0.312f

C12 IN1 GND 0.339f

C13 a_n12_34# GND 0.0101f **FLOATING

C14 a_n12_166# GND 0.671f **FLOATING

C15 w_n86_148# GND 1.33f **FLOATING

//.ends

.tran 1n 20n

.control

run

.endc

.end
