magic
tech sky130A
timestamp 1737132347
<< error_p >>
rect 93 103 94 121
<< nwell >>
rect -98 -15 442 143
<< nmos >>
rect -18 -141 -3 -99
rect 98 -141 113 -97
rect 148 -141 163 -97
rect 198 -141 213 -97
rect 248 -141 263 -97
rect 367 -141 382 -97
<< pmos >>
rect -18 9 -3 53
rect 98 9 113 53
rect 148 9 163 53
rect 198 9 213 53
rect 248 9 263 53
rect 367 9 382 54
<< ndiff >>
rect -53 -107 -18 -99
rect -53 -135 -43 -107
rect -26 -135 -18 -107
rect -53 -141 -18 -135
rect -3 -107 32 -99
rect -3 -135 6 -107
rect 23 -135 32 -107
rect -3 -141 32 -135
rect 64 -105 98 -97
rect 64 -133 72 -105
rect 89 -133 98 -105
rect 64 -141 98 -133
rect 113 -141 148 -97
rect 163 -105 198 -97
rect 163 -133 172 -105
rect 189 -133 198 -105
rect 163 -141 198 -133
rect 213 -141 248 -97
rect 263 -105 295 -97
rect 263 -133 271 -105
rect 288 -133 295 -105
rect 263 -141 295 -133
rect 333 -105 367 -97
rect 333 -133 343 -105
rect 360 -133 367 -105
rect 333 -141 367 -133
rect 382 -105 416 -97
rect 382 -133 392 -105
rect 409 -133 416 -105
rect 382 -141 416 -133
<< pdiff >>
rect -53 46 -18 53
rect -53 17 -45 46
rect -27 17 -18 46
rect -53 9 -18 17
rect -3 46 32 53
rect -3 17 6 46
rect 24 17 32 46
rect -3 9 32 17
rect 63 45 98 53
rect 63 16 71 45
rect 89 16 98 45
rect 63 9 98 16
rect 113 45 148 53
rect 113 16 122 45
rect 139 16 148 45
rect 113 9 148 16
rect 163 46 198 53
rect 163 17 172 46
rect 189 17 198 46
rect 163 9 198 17
rect 213 46 248 53
rect 213 17 222 46
rect 239 17 248 46
rect 213 9 248 17
rect 263 46 301 53
rect 263 17 274 46
rect 291 17 301 46
rect 263 9 301 17
rect 333 46 367 54
rect 333 17 342 46
rect 359 17 367 46
rect 333 9 367 17
rect 382 45 417 54
rect 382 16 392 45
rect 409 16 417 45
rect 382 9 417 16
<< ndiffc >>
rect -43 -135 -26 -107
rect 6 -135 23 -107
rect 72 -133 89 -105
rect 172 -133 189 -105
rect 271 -133 288 -105
rect 343 -133 360 -105
rect 392 -133 409 -105
<< pdiffc >>
rect -45 17 -27 46
rect 6 17 24 46
rect 71 16 89 45
rect 122 16 139 45
rect 172 17 189 46
rect 222 17 239 46
rect 274 17 291 46
rect 342 17 359 46
rect 392 16 409 45
<< psubdiff >>
rect -101 -173 442 -168
rect -101 -191 -10 -173
rect 7 -191 28 -173
rect 45 -191 108 -173
rect 125 -191 151 -173
rect 168 -191 194 -173
rect 211 -191 237 -173
rect 254 -191 305 -173
rect 322 -191 387 -173
rect 404 -191 442 -173
rect -101 -197 442 -191
<< nsubdiff >>
rect -72 122 424 125
rect -72 121 379 122
rect -72 119 24 121
rect -72 101 -12 119
rect 5 103 24 119
rect 41 120 93 121
rect 41 103 60 120
rect 5 102 60 103
rect 77 103 93 120
rect 110 103 162 121
rect 179 120 313 121
rect 179 103 200 120
rect 77 102 200 103
rect 217 119 276 120
rect 217 102 240 119
rect 5 101 240 102
rect 257 102 276 119
rect 293 103 313 120
rect 330 104 379 121
rect 396 104 424 122
rect 330 103 424 104
rect 293 102 424 103
rect 257 101 424 102
rect -72 96 424 101
<< psubdiffcont >>
rect -10 -191 7 -173
rect 28 -191 45 -173
rect 108 -191 125 -173
rect 151 -191 168 -173
rect 194 -191 211 -173
rect 237 -191 254 -173
rect 305 -191 322 -173
rect 387 -191 404 -173
<< nsubdiffcont >>
rect -12 101 5 119
rect 24 103 41 121
rect 60 102 77 120
rect 93 103 110 121
rect 162 103 179 121
rect 200 102 217 120
rect 240 101 257 119
rect 276 102 293 120
rect 313 103 330 121
rect 379 104 396 122
<< poly >>
rect -18 53 -3 75
rect 98 53 113 75
rect 148 53 163 75
rect 198 53 213 75
rect 248 53 263 75
rect 367 54 382 75
rect -18 -99 -3 9
rect 98 -97 113 9
rect 148 -97 163 9
rect 198 -12 213 9
rect 184 -20 213 -12
rect 184 -37 189 -20
rect 206 -37 213 -20
rect 184 -45 213 -37
rect 198 -97 213 -45
rect 248 -97 263 9
rect 313 -56 346 -49
rect 313 -73 321 -56
rect 338 -63 346 -56
rect 367 -63 382 9
rect 338 -73 382 -63
rect 313 -80 382 -73
rect 367 -97 382 -80
rect -18 -158 -3 -141
rect 98 -154 113 -141
rect 148 -154 163 -141
rect 198 -154 213 -141
rect 248 -154 263 -141
rect 367 -154 382 -141
<< polycont >>
rect 189 -37 206 -20
rect 321 -73 338 -56
<< locali >>
rect -95 122 442 125
rect -95 121 122 122
rect -95 119 24 121
rect -95 101 -82 119
rect -65 101 -46 119
rect -29 101 -12 119
rect 5 103 24 119
rect 41 120 93 121
rect 41 103 60 120
rect 5 102 60 103
rect 77 103 93 120
rect 110 104 122 121
rect 139 121 343 122
rect 139 104 162 121
rect 110 103 162 104
rect 179 120 313 121
rect 179 103 200 120
rect 77 102 200 103
rect 217 119 276 120
rect 217 102 240 119
rect 5 101 240 102
rect 257 102 276 119
rect 293 103 313 120
rect 330 104 343 121
rect 360 104 379 122
rect 396 104 442 122
rect 330 103 442 104
rect 293 102 442 103
rect 257 101 442 102
rect -95 96 442 101
rect -43 53 -26 96
rect 123 53 140 96
rect 344 54 361 96
rect -53 46 -19 53
rect -53 17 -45 46
rect -27 17 -19 46
rect -53 9 -19 17
rect -2 46 32 53
rect -2 17 6 46
rect 24 17 32 46
rect -2 9 32 17
rect 63 45 97 53
rect 63 16 71 45
rect 89 16 97 45
rect 63 9 97 16
rect 114 45 147 53
rect 114 16 122 45
rect 139 16 147 45
rect 114 9 147 16
rect 164 46 197 53
rect 164 17 172 46
rect 189 17 197 46
rect 164 9 197 17
rect 214 46 247 53
rect 214 17 222 46
rect 239 17 247 46
rect 214 9 247 17
rect 264 46 301 53
rect 264 17 274 46
rect 291 17 301 46
rect 264 9 301 17
rect 333 46 366 54
rect 333 17 342 46
rect 359 17 366 46
rect 333 9 366 17
rect 383 45 417 54
rect 383 16 392 45
rect 409 16 417 45
rect 383 9 417 16
rect 7 -20 24 9
rect 184 -20 213 -12
rect 7 -37 189 -20
rect 206 -37 213 -20
rect 7 -99 24 -37
rect 184 -45 213 -37
rect 230 -63 247 9
rect 395 -40 412 9
rect 313 -56 346 -49
rect 313 -63 321 -56
rect 171 -73 321 -63
rect 338 -73 346 -56
rect 171 -80 346 -73
rect 395 -57 439 -40
rect 171 -97 188 -80
rect 395 -97 412 -57
rect -53 -107 -19 -99
rect -53 -135 -43 -107
rect -26 -135 -19 -107
rect -53 -141 -19 -135
rect -2 -107 32 -99
rect -2 -135 6 -107
rect 23 -135 32 -107
rect -2 -141 32 -135
rect 64 -105 97 -97
rect 64 -133 72 -105
rect 89 -133 97 -105
rect 64 -141 97 -133
rect 164 -105 195 -97
rect 164 -133 172 -105
rect 189 -133 195 -105
rect 164 -141 195 -133
rect 264 -105 295 -97
rect 264 -133 271 -105
rect 288 -133 295 -105
rect 264 -141 295 -133
rect 333 -105 366 -97
rect 333 -133 343 -105
rect 360 -133 366 -105
rect 333 -141 366 -133
rect 383 -105 416 -97
rect 383 -133 392 -105
rect 409 -133 416 -105
rect 383 -141 416 -133
rect -43 -168 -26 -141
rect 71 -168 88 -141
rect 270 -168 287 -141
rect 343 -168 360 -141
rect -101 -173 442 -168
rect -101 -191 -83 -173
rect -66 -191 -42 -173
rect -25 -191 -10 -173
rect 7 -191 28 -173
rect 45 -191 71 -173
rect 88 -191 108 -173
rect 125 -191 151 -173
rect 168 -191 194 -173
rect 211 -191 237 -173
rect 254 -191 269 -173
rect 286 -191 305 -173
rect 322 -191 343 -173
rect 360 -191 387 -173
rect 404 -191 442 -173
rect -101 -197 442 -191
<< viali >>
rect -82 101 -65 119
rect -46 101 -29 119
rect 122 104 139 122
rect 343 104 360 122
rect 71 16 88 45
rect 172 17 189 46
rect 274 17 291 46
rect -83 -191 -66 -173
rect -42 -191 -25 -173
rect 71 -191 88 -173
rect 269 -191 286 -173
rect 343 -191 360 -173
<< metal1 >>
rect -95 122 442 125
rect -95 119 122 122
rect -95 101 -82 119
rect -65 101 -46 119
rect -29 104 122 119
rect 139 104 343 122
rect 360 104 442 122
rect -29 101 442 104
rect -95 96 442 101
rect 63 45 97 53
rect 63 16 71 45
rect 88 38 97 45
rect 164 46 197 53
rect 164 38 172 46
rect 88 20 172 38
rect 88 16 97 20
rect 63 9 97 16
rect 164 17 172 20
rect 189 38 197 46
rect 264 46 301 53
rect 264 38 274 46
rect 189 20 274 38
rect 189 17 197 20
rect 164 9 197 17
rect 264 17 274 20
rect 291 17 301 46
rect 264 9 301 17
rect -101 -173 442 -168
rect -101 -191 -83 -173
rect -66 -191 -42 -173
rect -25 -191 71 -173
rect 88 -191 269 -173
rect 286 -191 343 -173
rect 360 -191 442 -173
rect -101 -197 442 -191
<< labels >>
flabel metal1 s -87 102 -60 119 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel metal1 s -93 -190 -66 -173 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel poly s 247 -156 268 -140 0 FreeSans 80 0 0 0 I0
port 2 nsew
flabel poly s 97 -156 118 -140 0 FreeSans 80 0 0 0 I1
port 3 nsew
flabel poly s 146 -154 167 -138 0 FreeSans 80 0 0 0 S
port 4 nsew
flabel poly s -21 -159 0 -143 0 FreeSans 80 0 0 0 S
flabel locali s 410 -57 431 -41 0 FreeSans 80 0 0 0 OUT
port 5 nsew
<< end >>
