* SPICE3 file created from DFF.ext - technology: sky130A
.include pshort.lib
.include nshort.lib
.option scale=0.01u

//.subckt DFF VDD GND D CLK Q
M1000 a_606_n141# a_494_n141# GND GND nshort_model.0 ad=1470 pd=154 as=1470 ps=154 w=42 l=15
M1001 a_606_n141# a_494_n141# VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1002 a_772_n141# a_606_n141# a_672_9# VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1003 a_113_n141# D GND GND nshort_model.0 ad=770 pd=79u as=1500 ps=156 w=44 l=15
M1004 a_n3_n141# CLK VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1005 a_213_n141# a_n3_n141# a_163_n141# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1006 a_772_n141# a_494_n141# a_722_n141# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1007 a_163_n141# a_n3_n141# a_63_9# VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1008 Q a_772_n141# VDD VDD pshort_model.0 ad=1580 pd=160 as=1530 ps=158 w=45 l=15
M1009 Q a_772_n141# GND GND nshort_model.0 ad=1500 pd=156 as=1500 ps=156 w=44 l=15
M1010 a_63_9# CLK VDD VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1011 GND a_248_n154# a_213_n141# GND nshort_model.0 ad=1410 pd=152 as=770 ps=79u w=44 l=15
M1012 a_822_n141# a_606_n141# a_772_n141# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1013 VDD D a_63_9# VDD pshort_model.0 ad=770 pd=79u as=1540 ps=158 w=44 l=15
M1014 a_494_n141# CLK VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1015 a_63_9# a_248_n154# a_163_n141# VDD pshort_model.0 ad=1670 pd=164 as=770 ps=79u w=44 l=15
M1016 a_163_n141# CLK a_113_n141# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1017 a_722_n141# a_248_n154# GND GND nshort_model.0 ad=770 pd=79u as=1500 ps=156 w=44 l=15
M1018 a_672_9# a_494_n141# VDD VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1019 a_n3_n141# CLK GND GND nshort_model.0 ad=1470 pd=154 as=1470 ps=154 w=42 l=15
M1020 a_494_n141# CLK GND GND nshort_model.0 ad=1470 pd=154 as=1470 ps=154 w=42 l=15
M1021 a_248_n154# a_163_n141# GND GND nshort_model.0 ad=1500 pd=156 as=1500 ps=156 w=44 l=15
M1022 VDD a_248_n154# a_672_9# VDD pshort_model.0 ad=770 pd=79u as=1540 ps=158 w=44 l=15
M1023 a_672_9# Q a_772_n141# VDD pshort_model.0 ad=1670 pd=164 as=770 ps=79u w=44 l=15
M1024 GND Q a_822_n141# GND nshort_model.0 ad=1410 pd=152 as=770 ps=79u w=44 l=15
M1025 a_248_n154# a_163_n141# VDD VDD pshort_model.0 ad=1580 pd=160 as=1530 ps=158 w=45 l=15

VDD VDD 0 5V
VSS VSS 0 0V
Va D VSS PULSE(0 5V 0 0.1ns 0.1ns 3ns 9ns)
Vb CLK VSS PULSE(0 5V 0 0.1ns 0.1ns 2ns 4ns)

C0 a_n3_n141# a_163_n141# 0.15f
C1 a_672_9# a_494_n141# 0.0451f
C2 CLK a_113_n141# 0.00346f
C3 a_772_n141# a_722_n141# 0.00374f
C4 a_772_n141# VDD 0.0507f
C5 a_248_n154# CLK 0.212f
C6 a_248_n154# Q 6.5e-19
C7 a_248_n154# a_494_n141# 0.466f
C8 a_606_n141# a_672_9# 0.184f
C9 a_63_9# VDD 0.551f
C10 a_163_n141# a_113_n141# 0.00374f
C11 a_494_n141# CLK 0.146f
C12 a_494_n141# Q 7.72e-19
C13 a_163_n141# a_248_n154# 0.332f
C14 a_163_n141# CLK 0.159f
C15 a_n3_n141# VDD 0.219f
C16 a_672_9# a_722_n141# 5.89e-19
C17 a_672_9# VDD 0.55f
C18 a_163_n141# a_494_n141# 2.87e-19
C19 a_248_n154# a_606_n141# 0.133f
C20 a_606_n141# Q 0.0928f
C21 a_606_n141# a_494_n141# 0.315f
C22 a_248_n154# a_722_n141# 0.00157f
C23 a_248_n154# VDD 0.266f
C24 CLK VDD 0.177f
C25 Q VDD 0.197f
C26 a_63_9# D 0.0108f
C27 a_248_n154# a_213_n141# 0.00117f
C28 a_494_n141# a_722_n141# 0.00395f
C29 a_494_n141# VDD 0.256f
C30 a_213_n141# CLK 0.00197f
C31 a_n3_n141# D 0.0219f
C32 a_772_n141# a_822_n141# 0.00738f
C33 a_163_n141# VDD 0.0503f
C34 a_163_n141# a_213_n141# 0.00738f
C35 a_606_n141# a_722_n141# 0.00167f
C36 a_606_n141# VDD 0.202f
C37 D CLK 0.15f
C38 a_672_9# a_822_n141# 0.00137f
C39 a_772_n141# a_672_9# 0.211f
C40 a_163_n141# D 0.00275f
C41 a_n3_n141# a_63_9# 0.213f
C42 a_248_n154# a_822_n141# 0.0011f
C43 a_248_n154# a_772_n141# 0.00591f
C44 a_772_n141# Q 0.325f
C45 D VDD 0.0129f
C46 a_63_9# a_248_n154# 0.0928f
C47 a_772_n141# a_494_n141# 0.0649f
C48 a_63_9# CLK 0.158f
C49 a_n3_n141# a_113_n141# 0.00162f
C50 a_n3_n141# a_248_n154# 0.0932f
C51 a_n3_n141# CLK 0.319f
C52 a_63_9# a_494_n141# 1.36e-19
C53 a_248_n154# a_672_9# 0.0413f
C54 a_672_9# CLK 4.7e-19
C55 a_672_9# Q 0.0897f
C56 a_63_9# a_163_n141# 0.205f
C57 a_606_n141# a_772_n141# 0.163f
C58 Q GND 0.536f
C59 D GND 0.171f
C60 CLK GND 1.17f
C61 VDD GND 3.95f
//C62 a_822_n141# GND 0.00921f **FLOATING
//C63 a_722_n141# GND 0.00921f **FLOATING
//C64 a_213_n141# GND 0.00921f **FLOATING
//C65 a_113_n141# GND 0.00921f **FLOATING
//C66 a_672_9# GND 0.115f **FLOATING
//C67 a_772_n141# GND 0.602f **FLOATING
//C68 a_606_n141# GND 0.467f **FLOATING
//C69 a_494_n141# GND 0.981f **FLOATING
//C70 a_63_9# GND 0.0689f **FLOATING
//C71 a_163_n141# GND 0.573f **FLOATING
//C72 a_248_n154# GND 1.34f **FLOATING
//C73 a_n3_n141# GND 0.509f **FLOATING
//.ends
.tran 1n 20n
.control
run
.endc
.end
