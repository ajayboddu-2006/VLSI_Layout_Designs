magic

tech sky130A

timestamp 1738390936

<< nwell >>

rect -161 87 1265 309

rect -161 86 -8 87

<< nmos >>

rect -89 -128 -71 -48

rect 60 -127 78 -47

rect 228 -127 246 -47

rect 300 -127 318 -47

rect 446 -127 464 -47

rect 592 -127 610 -47

rect 664 -127 682 -47

rect 810 -127 828 -47

rect 958 -127 976 -47

rect 1030 -127 1048 -47

rect 1176 -127 1194 -47

<< pmos >>

rect -89 125 -71 202

rect 60 126 78 203

rect 228 127 246 203

rect 300 127 318 203

rect 446 126 464 203

rect 592 127 610 203

rect 664 127 682 203

rect 810 126 828 203

rect 958 127 976 203

rect 1030 127 1048 203

rect 1176 126 1194 203

<< ndiff >>

rect -139 -57 -89 -48

rect -139 -111 -126 -57

rect -102 -111 -89 -57

rect -139 -128 -89 -111

rect -71 -59 -21 -48

rect -71 -113 -55 -59

rect -31 -113 -21 -59

rect -71 -128 -21 -113

rect 10 -56 60 -47

rect 10 -110 23 -56

rect 47 -110 60 -56

rect 10 -127 60 -110

rect 78 -58 128 -47

rect 78 -112 94 -58

rect 118 -112 128 -58

rect 78 -127 128 -112

rect 177 -59 228 -47

rect 177 -113 191 -59

rect 216 -113 228 -59

rect 177 -127 228 -113

rect 246 -127 300 -47

rect 318 -58 369 -47

rect 318 -112 335 -58

rect 360 -112 369 -58

rect 318 -127 369 -112

rect 396 -56 446 -47

rect 396 -110 409 -56

rect 433 -110 446 -56

rect 396 -127 446 -110

rect 464 -58 514 -47

rect 464 -112 480 -58

rect 504 -112 514 -58

rect 464 -127 514 -112

rect 541 -59 592 -47

rect 541 -113 555 -59

rect 580 -113 592 -59

rect 541 -127 592 -113

rect 610 -57 664 -47

rect 610 -111 626 -57

rect 651 -111 664 -57

rect 610 -127 664 -111

rect 682 -58 733 -47

rect 682 -112 699 -58

rect 724 -112 733 -58

rect 682 -127 733 -112

rect 760 -56 810 -47

rect 760 -110 773 -56

rect 797 -110 810 -56

rect 760 -127 810 -110

rect 828 -58 878 -47

rect 828 -112 844 -58

rect 868 -112 878 -58

rect 828 -127 878 -112

rect 907 -59 958 -47

rect 907 -113 921 -59

rect 946 -113 958 -59

rect 907 -127 958 -113

rect 976 -57 1030 -47

rect 976 -111 992 -57

rect 1017 -111 1030 -57

rect 976 -127 1030 -111

rect 1048 -58 1099 -47

rect 1048 -112 1065 -58

rect 1090 -112 1099 -58

rect 1048 -127 1099 -112

rect 1126 -56 1176 -47

rect 1126 -110 1139 -56

rect 1163 -110 1176 -56

rect 1126 -127 1176 -110

rect 1194 -58 1244 -47

rect 1194 -112 1210 -58

rect 1234 -112 1244 -58

rect 1194 -127 1244 -112

<< pdiff >>

rect -141 193 -89 202

rect -141 136 -128 193

rect -98 136 -89 193

rect -141 125 -89 136

rect -71 192 -19 202

rect -71 135 -58 192

rect -28 135 -19 192

rect -71 125 -19 135

rect 8 194 60 203

rect 8 137 21 194

rect 51 137 60 194

rect 8 126 60 137

rect 78 193 130 203

rect 78 136 91 193

rect 121 136 130 193

rect 78 126 130 136

rect 179 192 228 203

rect 179 139 192 192

rect 219 139 228 192

rect 179 127 228 139

rect 246 193 300 203

rect 246 140 263 193

rect 290 140 300 193

rect 246 127 300 140

rect 318 192 367 203

rect 318 139 330 192

rect 357 139 367 192

rect 318 127 367 139

rect 394 194 446 203

rect 394 137 407 194

rect 437 137 446 194

rect 394 126 446 137

rect 464 193 516 203

rect 464 136 477 193

rect 507 136 516 193

rect 464 126 516 136

rect 543 192 592 203

rect 543 139 556 192

rect 583 139 592 192

rect 543 127 592 139

rect 610 127 664 203

rect 682 192 731 203

rect 682 139 694 192

rect 721 139 731 192

rect 682 127 731 139

rect 758 194 810 203

rect 758 137 771 194

rect 801 137 810 194

rect 758 126 810 137

rect 828 193 880 203

rect 828 136 841 193

rect 871 136 880 193

rect 828 126 880 136

rect 909 192 958 203

rect 909 139 922 192

rect 949 139 958 192

rect 909 127 958 139

rect 976 127 1030 203

rect 1048 192 1097 203

rect 1048 139 1060 192

rect 1087 139 1097 192

rect 1048 127 1097 139

rect 1124 194 1176 203

rect 1124 137 1137 194

rect 1167 137 1176 194

rect 1124 126 1176 137

rect 1194 193 1246 203

rect 1194 136 1207 193

rect 1237 136 1246 193

rect 1194 126 1246 136

<< ndiffc >>

rect -126 -111 -102 -57

rect -55 -113 -31 -59

rect 23 -110 47 -56

rect 94 -112 118 -58

rect 191 -113 216 -59

rect 335 -112 360 -58

rect 409 -110 433 -56

rect 480 -112 504 -58

rect 555 -113 580 -59

rect 626 -111 651 -57

rect 699 -112 724 -58

rect 773 -110 797 -56

rect 844 -112 868 -58

rect 921 -113 946 -59

rect 992 -111 1017 -57

rect 1065 -112 1090 -58

rect 1139 -110 1163 -56

rect 1210 -112 1234 -58

<< pdiffc >>

rect -128 136 -98 193

rect -58 135 -28 192

rect 21 137 51 194

rect 91 136 121 193

rect 192 139 219 192

rect 263 140 290 193

rect 330 139 357 192

rect 407 137 437 194

rect 477 136 507 193

rect 556 139 583 192

rect 694 139 721 192

rect 771 137 801 194

rect 841 136 871 193

rect 922 139 949 192

rect 1060 139 1087 192

rect 1137 137 1167 194

rect 1207 136 1237 193

<< psubdiff >>

rect -142 -181 1256 -175

rect -142 -182 264 -181

rect -142 -184 151 -182

rect -142 -186 -30 -184

rect -142 -206 -78 -186

rect -57 -204 -30 -186

rect -9 -204 52 -184

rect 73 -204 102 -184

rect 123 -202 151 -184

rect 172 -201 264 -182

rect 285 -201 305 -181

rect 326 -182 733 -181

rect 326 -201 359 -182

rect 172 -202 359 -201

rect 380 -184 600 -182

rect 380 -185 510 -184

rect 380 -202 452 -185

rect 123 -204 452 -202

rect -57 -205 452 -204

rect 473 -204 510 -185

rect 531 -202 600 -184

rect 621 -202 653 -182

rect 674 -201 733 -182

rect 754 -184 1256 -181

rect 754 -201 837 -184

rect 674 -202 837 -201

rect 531 -204 837 -202

rect 858 -204 893 -184

rect 914 -204 982 -184

rect 1003 -204 1027 -184

rect 1048 -204 1103 -184

rect 1124 -185 1256 -184

rect 1124 -204 1187 -185

rect 473 -205 1187 -204

rect 1208 -205 1256 -185

rect -57 -206 1256 -205

rect -142 -211 1256 -206

<< nsubdiff >>

rect -142 281 1237 285

rect -142 280 739 281

rect -142 279 605 280

rect -142 278 106 279

rect -142 258 -76 278

rect -55 276 106 278

rect -55 258 61 276

rect -142 256 61 258

rect 82 259 106 276

rect 127 277 449 279

rect 127 259 154 277

rect 82 257 154 259

rect 175 257 240 277

rect 261 257 286 277

rect 307 276 449 277

rect 307 257 369 276

rect 82 256 369 257

rect 390 259 449 276

rect 470 276 605 279

rect 470 259 501 276

rect 390 256 501 259

rect 522 260 605 276

rect 626 279 739 280

rect 626 260 653 279

rect 522 259 653 260

rect 674 274 739 279

rect 674 259 698 274

rect 522 256 698 259

rect -142 254 698 256

rect 719 261 739 274

rect 760 279 1109 281

rect 760 261 819 279

rect 719 259 819 261

rect 840 259 877 279

rect 898 277 1109 279

rect 898 259 971 277

rect 719 257 971 259

rect 992 276 1071 277

rect 992 257 1021 276

rect 719 256 1021 257

rect 1042 257 1071 276

rect 1092 261 1109 277

rect 1130 279 1237 281

rect 1130 261 1189 279

rect 1092 259 1189 261

rect 1210 259 1237 279

rect 1092 257 1237 259

rect 1042 256 1237 257

rect 719 254 1237 256

rect -142 249 1237 254

<< psubdiffcont >>

rect -78 -206 -57 -186

rect -30 -204 -9 -184

rect 52 -204 73 -184

rect 102 -204 123 -184

rect 151 -202 172 -182

rect 264 -201 285 -181

rect 305 -201 326 -181

rect 359 -202 380 -182

rect 452 -205 473 -185

rect 510 -204 531 -184

rect 600 -202 621 -182

rect 653 -202 674 -182

rect 733 -201 754 -181

rect 837 -204 858 -184

rect 893 -204 914 -184

rect 982 -204 1003 -184

rect 1027 -204 1048 -184

rect 1103 -204 1124 -184

rect 1187 -205 1208 -185

<< nsubdiffcont >>

rect -76 258 -55 278

rect 61 256 82 276

rect 106 259 127 279

rect 154 257 175 277

rect 240 257 261 277

rect 286 257 307 277

rect 369 256 390 276

rect 449 259 470 279

rect 501 256 522 276

rect 605 260 626 280

rect 653 259 674 279

rect 698 254 719 274

rect 739 261 760 281

rect 819 259 840 279

rect 877 259 898 279

rect 971 257 992 277

rect 1021 256 1042 276

rect 1071 257 1092 277

rect 1109 261 1130 281

rect 1189 259 1210 279

<< poly >>

rect -89 202 -71 231

rect 60 203 78 232

rect 228 203 246 231

rect 300 203 318 230

rect 446 203 464 232

rect 592 203 610 231

rect 664 203 682 230

rect 810 203 828 232

rect 958 203 976 231

rect 1030 203 1048 230

rect 1176 203 1194 232

rect -89 -48 -71 125

rect 60 3 78 126

rect 228 110 246 127

rect 208 102 246 110

rect 208 81 216 102

rect 237 81 246 102

rect 208 73 246 81

rect 30 -2 78 3

rect 30 -24 39 -2

rect 59 -24 78 -2

rect 30 -30 78 -24

rect 60 -47 78 -30

rect 228 -47 246 73

rect 300 -47 318 127

rect 446 103 464 126

rect 592 104 610 127

rect 420 94 464 103

rect 420 72 431 94

rect 455 72 464 94

rect 420 62 464 72

rect 573 94 610 104

rect 573 74 583 94

rect 602 74 610 94

rect 573 66 610 74

rect 446 -47 464 62

rect 592 -47 610 66

rect 664 63 682 127

rect 810 107 828 126

rect 792 99 828 107

rect 792 77 799 99

rect 819 77 828 99

rect 792 69 828 77

rect 664 51 712 63

rect 664 31 684 51

rect 706 31 712 51

rect 664 22 712 31

rect 664 -47 682 22

rect 810 -47 828 69

rect 958 65 976 127

rect 932 52 976 65

rect 932 32 942 52

rect 964 32 976 52

rect 932 24 976 32

rect 958 -47 976 24

rect 1030 12 1048 127

rect 1176 109 1194 126

rect 1156 101 1194 109

rect 1156 79 1166 101

rect 1186 79 1194 101

rect 1156 71 1194 79

rect 1030 1 1074 12

rect 1030 -19 1046 1

rect 1068 -19 1074 1

rect 1030 -28 1074 -19

rect 1030 -47 1048 -28

rect 1176 -47 1194 71

rect -89 -153 -71 -128

rect 60 -152 78 -127

rect 228 -153 246 -127

rect 300 -154 318 -127

rect 446 -152 464 -127

rect 592 -153 610 -127

rect 664 -154 682 -127

rect 810 -152 828 -127

rect 958 -153 976 -127

rect 1030 -154 1048 -127

rect 1176 -152 1194 -127

<< polycont >>

rect 216 81 237 102

rect 39 -24 59 -2

rect 431 72 455 94

rect 583 74 602 94

rect 799 77 819 99

rect 684 31 706 51

rect 942 32 964 52

rect 1166 79 1186 101

rect 1046 -19 1068 1

<< locali >>

rect -142 281 1256 285

rect -142 280 739 281

rect -142 279 605 280

rect -142 278 106 279

rect -142 276 -76 278

rect -142 256 -126 276

rect -105 258 -76 276

rect -55 277 106 278

rect -55 258 23 277

rect -105 257 23 258

rect 44 276 106 277

rect 44 257 61 276

rect -105 256 61 257

rect 82 259 106 276

rect 127 277 449 279

rect 127 259 154 277

rect 82 257 154 259

rect 175 257 194 277

rect 215 257 240 277

rect 261 257 286 277

rect 307 276 409 277

rect 307 257 330 276

rect 82 256 330 257

rect 351 256 369 276

rect 390 257 409 276

rect 430 259 449 277

rect 470 277 605 279

rect 470 276 560 277

rect 470 259 501 276

rect 430 257 501 259

rect 390 256 501 257

rect 522 257 560 276

rect 581 260 605 277

rect 626 279 739 280

rect 626 260 653 279

rect 581 259 653 260

rect 674 274 739 279

rect 674 259 698 274

rect 581 257 698 259

rect 522 256 698 257

rect -142 254 698 256

rect 719 261 739 274

rect 760 279 1109 281

rect 760 277 819 279

rect 760 261 773 277

rect 719 257 773 261

rect 794 259 819 277

rect 840 259 877 279

rect 898 277 1109 279

rect 898 276 971 277

rect 898 259 926 276

rect 794 257 926 259

rect 719 256 926 257

rect 947 257 971 276

rect 992 276 1071 277

rect 992 257 1021 276

rect 947 256 1021 257

rect 1042 257 1071 276

rect 1092 261 1109 277

rect 1130 279 1256 281

rect 1130 277 1189 279

rect 1130 261 1139 277

rect 1092 257 1139 261

rect 1160 259 1189 277

rect 1210 259 1256 279

rect 1160 257 1256 259

rect 1042 256 1256 257

rect 719 254 1256 256

rect -142 249 1256 254

rect -126 202 -105 249

rect 23 203 44 249

rect 195 203 218 249

rect 331 246 359 249

rect 331 204 348 246

rect 331 203 359 204

rect 409 203 430 249

rect 559 203 582 249

rect 773 203 794 249

rect 925 203 948 249

rect 1139 203 1160 249

rect -141 193 -91 202

rect -141 136 -128 193

rect -98 136 -91 193

rect -141 125 -91 136

rect -69 192 -19 202

rect -69 135 -58 192

rect -28 135 -19 192

rect -69 125 -19 135

rect 8 194 58 203

rect 8 137 21 194

rect 51 137 58 194

rect 8 126 58 137

rect 80 193 130 203

rect 80 136 91 193

rect 121 136 130 193

rect 80 126 130 136

rect 179 192 226 203

rect 179 139 192 192

rect 219 139 226 192

rect 179 127 226 139

rect 249 193 296 203

rect 249 140 263 193

rect 290 140 296 193

rect 249 127 296 140

rect 320 192 367 203

rect 320 139 330 192

rect 357 139 367 192

rect 320 127 367 139

rect 394 194 444 203

rect 394 137 407 194

rect 437 137 444 194

rect -55 -48 -34 125

rect 94 97 115 126

rect 208 102 244 110

rect 208 97 216 102

rect 94 81 216 97

rect 237 81 244 102

rect 262 103 285 127

rect 394 126 444 137

rect 466 193 516 203

rect 466 136 477 193

rect 507 136 516 193

rect 466 126 516 136

rect 543 192 590 203

rect 543 139 556 192

rect 583 139 590 192

rect 543 127 590 139

rect 684 192 731 203

rect 684 139 694 192

rect 721 139 731 192

rect 684 127 731 139

rect 758 194 808 203

rect 758 137 771 194

rect 801 137 808 194

rect 262 94 463 103

rect 262 86 431 94

rect 94 80 244 81

rect 30 -2 67 3

rect 30 -24 39 -2

rect 59 -24 67 -2

rect 30 -30 67 -24

rect 94 -47 115 80

rect 208 73 244 80

rect 338 -47 359 86

rect 420 72 431 86

rect 455 72 463 94

rect 420 62 463 72

rect 480 99 501 126

rect 702 107 722 127

rect 758 126 808 137

rect 830 193 880 203

rect 830 136 841 193

rect 871 136 880 193

rect 830 126 880 136

rect 909 192 956 203

rect 909 139 922 192

rect 949 139 956 192

rect 909 127 956 139

rect 1050 192 1097 203

rect 1050 139 1060 192

rect 1087 139 1097 192

rect 1050 127 1097 139

rect 1124 194 1174 203

rect 1124 137 1137 194

rect 1167 137 1174 194

rect 573 99 609 104

rect 480 94 609 99

rect 480 79 583 94

rect 480 -47 501 79

rect 573 74 583 79

rect 602 74 609 94

rect 573 66 609 74

rect 629 99 826 107

rect 629 90 799 99

rect 629 -47 650 90

rect 792 77 799 90

rect 819 77 826 99

rect 792 69 826 77

rect 674 51 712 63

rect 674 31 684 51

rect 706 31 712 51

rect 674 22 712 31

rect 844 -47 865 126

rect 1072 103 1093 127

rect 1124 126 1174 137

rect 1196 193 1246 203

rect 1196 136 1207 193

rect 1237 136 1246 193

rect 1196 126 1246 136

rect 1156 103 1193 109

rect 992 101 1193 103

rect 992 85 1166 101

rect 932 52 970 65

rect 932 32 942 52

rect 964 32 970 52

rect 932 24 970 32

rect 992 -47 1014 85

rect 1156 79 1166 85

rect 1186 79 1193 101

rect 1156 71 1193 79

rect 1036 1 1074 12

rect 1036 -19 1046 1

rect 1068 -19 1074 1

rect 1036 -28 1074 -19

rect 1210 -47 1231 126

rect -139 -57 -91 -48

rect -139 -111 -126 -57

rect -102 -111 -91 -57

rect -139 -128 -91 -111

rect -69 -59 -21 -48

rect -69 -113 -55 -59

rect -31 -113 -21 -59

rect -69 -128 -21 -113

rect 10 -56 58 -47

rect 10 -110 23 -56

rect 47 -110 58 -56

rect 10 -127 58 -110

rect 80 -58 128 -47

rect 80 -112 94 -58

rect 118 -112 128 -58

rect 80 -127 128 -112

rect 177 -59 226 -47

rect 177 -113 191 -59

rect 216 -113 226 -59

rect 177 -127 226 -113

rect 320 -58 369 -47

rect 320 -112 335 -58

rect 360 -112 369 -58

rect 320 -127 369 -112

rect 396 -56 444 -47

rect 396 -110 409 -56

rect 433 -110 444 -56

rect 396 -127 444 -110

rect 466 -58 514 -47

rect 466 -112 480 -58

rect 504 -112 514 -58

rect 466 -127 514 -112

rect 541 -59 590 -47

rect 541 -113 555 -59

rect 580 -113 590 -59

rect 541 -127 590 -113

rect 612 -57 661 -47

rect 612 -111 626 -57

rect 651 -111 661 -57

rect 612 -127 661 -111

rect 684 -58 733 -47

rect 684 -112 699 -58

rect 724 -112 733 -58

rect 684 -127 733 -112

rect 760 -56 808 -47

rect 760 -110 773 -56

rect 797 -110 808 -56

rect 760 -127 808 -110

rect 830 -58 878 -47

rect 830 -112 844 -58

rect 868 -112 878 -58

rect 830 -127 878 -112

rect 907 -59 956 -47

rect 907 -113 921 -59

rect 946 -113 956 -59

rect 907 -127 956 -113

rect 978 -57 1027 -47

rect 978 -111 992 -57

rect 1017 -111 1027 -57

rect 978 -127 1027 -111

rect 1050 -58 1099 -47

rect 1050 -112 1065 -58

rect 1090 -112 1099 -58

rect 1050 -127 1099 -112

rect 1126 -56 1174 -47

rect 1126 -110 1139 -56

rect 1163 -110 1174 -56

rect 1126 -127 1174 -110

rect 1196 -58 1244 -47

rect 1196 -112 1210 -58

rect 1234 -112 1244 -58

rect 1196 -127 1244 -112

rect -126 -175 -107 -128

rect 23 -175 42 -127

rect 190 -175 213 -127

rect 409 -175 428 -127

rect 554 -175 577 -127

rect 699 -175 722 -127

rect 773 -175 792 -127

rect 920 -175 943 -127

rect 1065 -175 1088 -127

rect 1139 -175 1158 -127

rect -142 -180 1256 -175

rect -142 -181 694 -180

rect -142 -182 264 -181

rect -142 -183 22 -182

rect -142 -203 -123 -183

rect -102 -184 22 -183

rect -102 -186 -30 -184

rect -102 -203 -78 -186

rect -142 -206 -78 -203

rect -57 -204 -30 -186

rect -9 -202 22 -184

rect 43 -184 151 -182

rect 43 -202 52 -184

rect -9 -204 52 -202

rect 73 -204 102 -184

rect 123 -202 151 -184

rect 172 -183 264 -182

rect 172 -202 189 -183

rect 123 -203 189 -202

rect 210 -201 264 -183

rect 285 -201 305 -181

rect 326 -182 552 -181

rect 326 -201 359 -182

rect 210 -202 359 -201

rect 380 -183 552 -182

rect 380 -202 409 -183

rect 210 -203 409 -202

rect 430 -184 552 -183

rect 430 -185 510 -184

rect 430 -203 452 -185

rect 123 -204 452 -203

rect -57 -205 452 -204

rect 473 -204 510 -185

rect 531 -201 552 -184

rect 573 -182 694 -181

rect 573 -201 600 -182

rect 531 -202 600 -201

rect 621 -202 653 -182

rect 674 -200 694 -182

rect 715 -181 1256 -180

rect 715 -200 733 -181

rect 674 -201 733 -200

rect 754 -182 1256 -181

rect 754 -201 774 -182

rect 674 -202 774 -201

rect 795 -184 920 -182

rect 795 -202 837 -184

rect 531 -204 837 -202

rect 858 -204 893 -184

rect 914 -202 920 -184

rect 941 -184 1063 -182

rect 941 -202 982 -184

rect 914 -204 982 -202

rect 1003 -204 1027 -184

rect 1048 -202 1063 -184

rect 1084 -184 1142 -182

rect 1084 -202 1103 -184

rect 1048 -204 1103 -202

rect 1124 -202 1142 -184

rect 1163 -185 1256 -182

rect 1163 -202 1187 -185

rect 1124 -204 1187 -202

rect 473 -205 1187 -204

rect 1208 -205 1256 -185

rect -57 -206 1256 -205

rect -142 -211 1256 -206

<< viali >>

rect -126 256 -105 276

rect 23 257 44 277

rect 194 257 215 277

rect 330 256 351 276

rect 409 257 430 277

rect 560 257 581 277

rect 773 257 794 277

rect 926 256 947 276

rect 1139 257 1160 277

rect 39 -24 59 -2

rect 684 31 706 51

rect 942 32 964 52

rect 1046 -19 1068 1

rect -123 -203 -102 -183

rect 22 -202 43 -182

rect 189 -203 210 -183

rect 409 -203 430 -183

rect 552 -201 573 -181

rect 694 -200 715 -180

rect 774 -202 795 -182

rect 920 -202 941 -182

rect 1063 -202 1084 -182

rect 1142 -202 1163 -182

<< metal1 >>

rect -142 277 1256 285

rect -142 276 23 277

rect -142 256 -126 276

rect -105 257 23 276

rect 44 257 194 277

rect 215 276 409 277

rect 215 257 330 276

rect -105 256 330 257

rect 351 257 409 276

rect 430 257 560 277

rect 581 257 773 277

rect 794 276 1139 277

rect 794 257 926 276

rect 351 256 926 257

rect 947 257 1139 276

rect 1160 257 1256 277

rect 947 256 1256 257

rect -142 249 1256 256

rect 674 54 712 63

rect 932 54 976 65

rect 674 52 976 54

rect 674 51 942 52

rect 674 31 684 51

rect 706 35 942 51

rect 706 31 712 35

rect 674 22 712 31

rect 932 32 942 35

rect 964 32 976 52

rect 932 24 976 32

rect 30 -2 67 3

rect 30 -24 39 -2

rect 59 -6 67 -2

rect 1036 1 1074 12

rect 1036 -6 1046 1

rect 59 -19 1046 -6

rect 1068 -19 1074 1

rect 59 -23 1074 -19

rect 59 -24 67 -23

rect 30 -30 67 -24

rect 1036 -28 1074 -23

rect -142 -180 1256 -175

rect -142 -181 694 -180

rect -142 -182 552 -181

rect -142 -183 22 -182

rect -142 -203 -123 -183

rect -102 -202 22 -183

rect 43 -183 552 -182

rect 43 -202 189 -183

rect -102 -203 189 -202

rect 210 -203 409 -183

rect 430 -201 552 -183

rect 573 -200 694 -181

rect 715 -182 1256 -180

rect 715 -200 774 -182

rect 573 -201 774 -200

rect 430 -202 774 -201

rect 795 -202 920 -182

rect 941 -202 1063 -182

rect 1084 -202 1142 -182

rect 1163 -202 1256 -182

rect 430 -203 1256 -202

rect -142 -211 1256 -203

<< labels >>

flabel locali s -35 249 21 279 0 FreeSans 80 0 0 0 VDD

port 0 nsew

flabel locali s -24 -211 32 -181 0 FreeSans 80 0 0 0 GND

port 1 nsew

flabel poly s -99 -160 -58 -134 0 FreeSans 80 0 0 0 I0

port 2 nsew

flabel poly s 291 -158 332 -132 0 FreeSans 80 0 0 0 I1

port 3 nsew

flabel poly s 50 -157 91 -131 0 FreeSans 80 0 0 0 I2

port 4 nsew

flabel poly s 651 -160 692 -134 0 FreeSans 80 0 0 0 I3

port 5 nsew

flabel locali s 844 0 885 26 0 FreeSans 80 0 0 0 O0

port 6 nsew

flabel locali s 1206 22 1247 48 0 FreeSans 80 0 0 0 O1

port 7 nsew

<< end >>
