magic

tech sky130A

timestamp 1738331326

<< nwell >>

rect -98 -15 1051 143

<< nmos >>

rect -18 -141 -3 -99

rect 98 -141 113 -97

rect 148 -141 163 -97

rect 198 -141 213 -97

rect 248 -141 263 -97

rect 367 -141 382 -97

rect 479 -141 494 -99

rect 591 -141 606 -99

rect 707 -141 722 -97

rect 757 -141 772 -97

rect 807 -141 822 -97

rect 857 -141 872 -97

rect 976 -141 991 -97

<< pmos >>

rect -18 9 -3 53

rect 98 9 113 53

rect 148 9 163 53

rect 198 9 213 53

rect 248 9 263 53

rect 367 9 382 54

rect 479 9 494 53

rect 591 9 606 53

rect 707 9 722 53

rect 757 9 772 53

rect 807 9 822 53

rect 857 9 872 53

rect 976 9 991 54

<< ndiff >>

rect -53 -107 -18 -99

rect -53 -135 -43 -107

rect -26 -135 -18 -107

rect -53 -141 -18 -135

rect -3 -107 32 -99

rect -3 -135 6 -107

rect 23 -135 32 -107

rect -3 -141 32 -135

rect 64 -105 98 -97

rect 64 -133 72 -105

rect 89 -133 98 -105

rect 64 -141 98 -133

rect 113 -141 148 -97

rect 163 -105 198 -97

rect 163 -133 172 -105

rect 189 -133 198 -105

rect 163 -141 198 -133

rect 213 -141 248 -97

rect 263 -105 295 -97

rect 263 -133 271 -105

rect 288 -133 295 -105

rect 263 -141 295 -133

rect 333 -105 367 -97

rect 333 -133 343 -105

rect 360 -133 367 -105

rect 333 -141 367 -133

rect 382 -105 416 -97

rect 382 -133 392 -105

rect 409 -133 416 -105

rect 382 -141 416 -133

rect 444 -107 479 -99

rect 444 -135 454 -107

rect 471 -135 479 -107

rect 444 -141 479 -135

rect 494 -107 529 -99

rect 494 -135 503 -107

rect 520 -135 529 -107

rect 494 -141 529 -135

rect 556 -107 591 -99

rect 556 -135 566 -107

rect 583 -135 591 -107

rect 556 -141 591 -135

rect 606 -107 641 -99

rect 606 -135 615 -107

rect 632 -135 641 -107

rect 606 -141 641 -135

rect 673 -105 707 -97

rect 673 -133 681 -105

rect 698 -133 707 -105

rect 673 -141 707 -133

rect 722 -141 757 -97

rect 772 -105 807 -97

rect 772 -133 781 -105

rect 798 -133 807 -105

rect 772 -141 807 -133

rect 822 -141 857 -97

rect 872 -105 904 -97

rect 872 -133 880 -105

rect 897 -133 904 -105

rect 872 -141 904 -133

rect 942 -105 976 -97

rect 942 -133 952 -105

rect 969 -133 976 -105

rect 942 -141 976 -133

rect 991 -105 1025 -97

rect 991 -133 1001 -105

rect 1018 -133 1025 -105

rect 991 -141 1025 -133

<< pdiff >>

rect -53 46 -18 53

rect -53 17 -45 46

rect -27 17 -18 46

rect -53 9 -18 17

rect -3 46 32 53

rect -3 17 6 46

rect 24 17 32 46

rect -3 9 32 17

rect 63 45 98 53

rect 63 16 71 45

rect 89 16 98 45

rect 63 9 98 16

rect 113 45 148 53

rect 113 16 122 45

rect 139 16 148 45

rect 113 9 148 16

rect 163 46 198 53

rect 163 17 172 46

rect 189 17 198 46

rect 163 9 198 17

rect 213 46 248 53

rect 213 17 222 46

rect 239 17 248 46

rect 213 9 248 17

rect 263 46 301 53

rect 263 17 274 46

rect 291 17 301 46

rect 263 9 301 17

rect 333 46 367 54

rect 333 17 342 46

rect 359 17 367 46

rect 333 9 367 17

rect 382 45 417 54

rect 382 16 392 45

rect 409 16 417 45

rect 382 9 417 16

rect 444 46 479 53

rect 444 17 452 46

rect 470 17 479 46

rect 444 9 479 17

rect 494 46 529 53

rect 494 17 503 46

rect 521 17 529 46

rect 494 9 529 17

rect 556 46 591 53

rect 556 17 564 46

rect 582 17 591 46

rect 556 9 591 17

rect 606 46 641 53

rect 606 17 615 46

rect 633 17 641 46

rect 606 9 641 17

rect 672 45 707 53

rect 672 16 680 45

rect 698 16 707 45

rect 672 9 707 16

rect 722 45 757 53

rect 722 16 731 45

rect 748 16 757 45

rect 722 9 757 16

rect 772 46 807 53

rect 772 17 781 46

rect 798 17 807 46

rect 772 9 807 17

rect 822 46 857 53

rect 822 17 831 46

rect 848 17 857 46

rect 822 9 857 17

rect 872 46 910 53

rect 872 17 883 46

rect 900 17 910 46

rect 872 9 910 17

rect 942 46 976 54

rect 942 17 951 46

rect 968 17 976 46

rect 942 9 976 17

rect 991 45 1026 54

rect 991 16 1001 45

rect 1018 16 1026 45

rect 991 9 1026 16

<< ndiffc >>

rect -43 -135 -26 -107

rect 6 -135 23 -107

rect 72 -133 89 -105

rect 172 -133 189 -105

rect 271 -133 288 -105

rect 343 -133 360 -105

rect 392 -133 409 -105

rect 454 -135 471 -107

rect 503 -135 520 -107

rect 566 -135 583 -107

rect 615 -135 632 -107

rect 681 -133 698 -105

rect 781 -133 798 -105

rect 880 -133 897 -105

rect 952 -133 969 -105

rect 1001 -133 1018 -105

<< pdiffc >>

rect -45 17 -27 46

rect 6 17 24 46

rect 71 16 89 45

rect 122 16 139 45

rect 172 17 189 46

rect 222 17 239 46

rect 274 17 291 46

rect 342 17 359 46

rect 392 16 409 45

rect 452 17 470 46

rect 503 17 521 46

rect 564 17 582 46

rect 615 17 633 46

rect 680 16 698 45

rect 731 16 748 45

rect 781 17 798 46

rect 831 17 848 46

rect 883 17 900 46

rect 951 17 968 46

rect 1001 16 1018 45

<< psubdiff >>

rect -101 -173 1051 -168

rect -101 -191 -10 -173

rect 7 -191 28 -173

rect 45 -191 108 -173

rect 125 -191 151 -173

rect 168 -191 194 -173

rect 211 -191 237 -173

rect 254 -191 305 -173

rect 322 -191 373 -173

rect 390 -191 487 -173

rect 504 -191 525 -173

rect 542 -191 599 -173

rect 616 -191 637 -173

rect 654 -191 717 -173

rect 734 -191 760 -173

rect 777 -191 803 -173

rect 820 -191 846 -173

rect 863 -191 914 -173

rect 931 -191 996 -173

rect 1013 -191 1051 -173

rect -101 -197 1051 -191

<< nsubdiff >>

rect -72 122 1033 125

rect -72 121 988 122

rect -72 119 24 121

rect -72 101 -12 119

rect 5 103 24 119

rect 41 120 94 121

rect 41 103 60 120

rect 5 102 60 103

rect 77 103 94 120

rect 111 103 162 121

rect 179 120 313 121

rect 179 103 200 120

rect 77 102 200 103

rect 217 119 276 120

rect 217 102 240 119

rect 5 101 240 102

rect 257 102 276 119

rect 293 103 313 120

rect 330 120 521 121

rect 330 103 374 120

rect 293 102 374 103

rect 391 119 521 120

rect 391 102 485 119

rect 257 101 485 102

rect 502 103 521 119

rect 538 119 633 121

rect 538 103 597 119

rect 502 101 597 103

rect 614 103 633 119

rect 650 120 703 121

rect 650 103 669 120

rect 614 102 669 103

rect 686 103 703 120

rect 720 103 771 121

rect 788 120 922 121

rect 788 103 809 120

rect 686 102 809 103

rect 826 119 885 120

rect 826 102 849 119

rect 614 101 849 102

rect 866 102 885 119

rect 902 103 922 120

rect 939 104 988 121

rect 1005 104 1033 122

rect 939 103 1033 104

rect 902 102 1033 103

rect 866 101 1033 102

rect -72 96 1033 101

<< psubdiffcont >>

rect -10 -191 7 -173

rect 28 -191 45 -173

rect 108 -191 125 -173

rect 151 -191 168 -173

rect 194 -191 211 -173

rect 237 -191 254 -173

rect 305 -191 322 -173

rect 373 -191 390 -173

rect 487 -191 504 -173

rect 525 -191 542 -173

rect 599 -191 616 -173

rect 637 -191 654 -173

rect 717 -191 734 -173

rect 760 -191 777 -173

rect 803 -191 820 -173

rect 846 -191 863 -173

rect 914 -191 931 -173

rect 996 -191 1013 -173

<< nsubdiffcont >>

rect -12 101 5 119

rect 24 103 41 121

rect 60 102 77 120

rect 94 103 111 121

rect 162 103 179 121

rect 200 102 217 120

rect 240 101 257 119

rect 276 102 293 120

rect 313 103 330 121

rect 374 102 391 120

rect 485 101 502 119

rect 521 103 538 121

rect 597 101 614 119

rect 633 103 650 121

rect 669 102 686 120

rect 703 103 720 121

rect 771 103 788 121

rect 809 102 826 120

rect 849 101 866 119

rect 885 102 902 120

rect 922 103 939 121

rect 988 104 1005 122

<< poly >>

rect -18 53 -3 75

rect 98 53 113 75

rect 148 53 163 75

rect 198 53 213 75

rect 248 53 263 75

rect 367 54 382 75

rect 479 53 494 75

rect 591 53 606 75

rect 707 53 722 75

rect 757 53 772 75

rect 807 53 822 75

rect 857 53 872 75

rect 976 54 991 75

rect -18 -51 -3 9

rect -43 -58 -3 -51

rect -43 -75 -35 -58

rect -18 -75 -3 -58

rect -43 -82 -3 -75

rect -42 -84 -3 -82

rect -18 -99 -3 -84

rect 98 -97 113 9

rect 148 -46 163 9

rect 198 -8 213 9

rect 184 -16 213 -8

rect 184 -33 189 -16

rect 206 -33 213 -16

rect 184 -45 213 -33

rect 134 -55 163 -46

rect 134 -72 141 -55

rect 158 -72 163 -55

rect 134 -80 163 -72

rect 148 -97 163 -80

rect 198 -97 213 -45

rect 248 -6 263 9

rect 248 -15 292 -6

rect 248 -32 269 -15

rect 286 -32 292 -15

rect 248 -40 292 -32

rect 248 -97 263 -40

rect 313 -56 346 -49

rect 313 -73 321 -56

rect 338 -63 346 -56

rect 367 -63 382 9

rect 479 -48 494 9

rect 338 -73 382 -63

rect 313 -80 382 -73

rect 453 -56 494 -48

rect 591 -49 606 9

rect 707 -47 722 9

rect 757 -47 772 9

rect 807 -12 822 9

rect 793 -20 822 -12

rect 793 -37 798 -20

rect 815 -37 822 -20

rect 793 -45 822 -37

rect 453 -73 461 -56

rect 478 -73 494 -56

rect 453 -80 494 -73

rect 367 -97 382 -80

rect 479 -99 494 -80

rect 566 -57 606 -49

rect 566 -74 574 -57

rect 591 -74 606 -57

rect 566 -81 606 -74

rect 591 -99 606 -81

rect 688 -56 722 -47

rect 688 -73 694 -56

rect 711 -73 722 -56

rect 688 -82 722 -73

rect 743 -55 772 -47

rect 743 -72 748 -55

rect 765 -72 772 -55

rect 743 -80 772 -72

rect 707 -97 722 -82

rect 757 -97 772 -80

rect 807 -97 822 -45

rect 857 -8 872 9

rect 857 -16 901 -8

rect 857 -33 879 -16

rect 896 -33 901 -16

rect 857 -41 901 -33

rect 857 -97 872 -41

rect 922 -56 955 -49

rect 922 -73 930 -56

rect 947 -63 955 -56

rect 976 -63 991 9

rect 947 -73 991 -63

rect 922 -80 991 -73

rect 976 -97 991 -80

rect -18 -158 -3 -141

rect 98 -154 113 -141

rect 148 -154 163 -141

rect 198 -154 213 -141

rect 248 -154 263 -141

rect 367 -154 382 -141

rect 479 -158 494 -141

rect 591 -158 606 -141

rect 707 -154 722 -141

rect 757 -154 772 -141

rect 807 -154 822 -141

rect 857 -154 872 -141

rect 976 -154 991 -141

<< polycont >>

rect -35 -75 -18 -58

rect 189 -33 206 -16

rect 141 -72 158 -55

rect 269 -32 286 -15

rect 321 -73 338 -56

rect 798 -37 815 -20

rect 461 -73 478 -56

rect 574 -74 591 -57

rect 694 -73 711 -56

rect 748 -72 765 -55

rect 879 -33 896 -16

rect 930 -73 947 -56

<< locali >>

rect -95 122 1051 125

rect -95 121 122 122

rect -95 119 24 121

rect -95 101 -82 119

rect -65 101 -46 119

rect -29 101 -12 119

rect 5 103 24 119

rect 41 120 94 121

rect 41 103 60 120

rect 5 102 60 103

rect 77 103 94 120

rect 111 104 122 121

rect 139 121 343 122

rect 139 104 162 121

rect 111 103 162 104

rect 179 120 313 121

rect 179 103 200 120

rect 77 102 200 103

rect 217 119 276 120

rect 217 102 240 119

rect 5 101 240 102

rect 257 102 276 119

rect 293 103 313 120

rect 330 104 343 121

rect 360 121 731 122

rect 360 120 521 121

rect 360 104 374 120

rect 330 103 374 104

rect 293 102 374 103

rect 391 119 521 120

rect 391 102 415 119

rect 257 101 415 102

rect 432 101 451 119

rect 468 101 485 119

rect 502 103 521 119

rect 538 119 633 121

rect 538 103 563 119

rect 502 101 563 103

rect 580 101 597 119

rect 614 103 633 119

rect 650 120 703 121

rect 650 103 669 120

rect 614 102 669 103

rect 686 103 703 120

rect 720 104 731 121

rect 748 121 952 122

rect 748 104 771 121

rect 720 103 771 104

rect 788 120 922 121

rect 788 103 809 120

rect 686 102 809 103

rect 826 119 885 120

rect 826 102 849 119

rect 614 101 849 102

rect 866 102 885 119

rect 902 103 922 120

rect 939 104 952 121

rect 969 104 988 122

rect 1005 104 1051 122

rect 939 103 1051 104

rect 902 102 1051 103

rect 866 101 1051 102

rect -95 96 1051 101

rect -43 53 -26 96

rect 123 53 140 96

rect 344 54 361 96

rect -53 46 -19 53

rect -53 17 -45 46

rect -27 17 -19 46

rect -53 9 -19 17

rect -2 46 32 53

rect -2 17 6 46

rect 24 17 32 46

rect -2 9 32 17

rect 63 45 97 53

rect 63 16 71 45

rect 89 16 97 45

rect 63 9 97 16

rect 114 45 147 53

rect 114 16 122 45

rect 139 16 147 45

rect 114 9 147 16

rect 164 46 197 53

rect 164 17 172 46

rect 189 17 197 46

rect 164 9 197 17

rect 214 46 247 53

rect 214 17 222 46

rect 239 17 247 46

rect 214 9 247 17

rect 264 46 301 53

rect 264 17 274 46

rect 291 17 301 46

rect 264 9 301 17

rect 333 46 366 54

rect 333 17 342 46

rect 359 17 366 46

rect 333 9 366 17

rect 383 45 417 54

rect 454 53 471 96

rect 566 53 583 96

rect 732 53 749 96

rect 953 54 970 96

rect 383 16 392 45

rect 409 16 417 45

rect 383 9 417 16

rect 444 46 478 53

rect 444 17 452 46

rect 470 17 478 46

rect 444 9 478 17

rect 495 46 529 53

rect 495 17 503 46

rect 521 17 529 46

rect 495 9 529 17

rect 556 46 590 53

rect 556 17 564 46

rect 582 17 590 46

rect 556 9 590 17

rect 607 46 641 53

rect 607 17 615 46

rect 633 17 641 46

rect 607 9 641 17

rect 672 45 706 53

rect 672 16 680 45

rect 698 16 706 45

rect 672 9 706 16

rect 723 45 756 53

rect 723 16 731 45

rect 748 16 756 45

rect 723 9 756 16

rect 773 46 806 53

rect 773 17 781 46

rect 798 17 806 46

rect 773 9 806 17

rect 823 46 856 53

rect 823 17 831 46

rect 848 17 856 46

rect 823 9 856 17

rect 873 46 910 53

rect 873 17 883 46

rect 900 17 910 46

rect 873 9 910 17

rect 942 46 975 54

rect 942 17 951 46

rect 968 17 975 46

rect 942 9 975 17

rect 992 45 1026 54

rect 992 16 1001 45

rect 1018 16 1026 45

rect 992 9 1026 16

rect 7 -8 24 9

rect 7 -16 210 -8

rect 7 -25 189 -16

rect -42 -51 -10 -50

rect -43 -58 -10 -51

rect -43 -75 -38 -58

rect -18 -75 -10 -58

rect -43 -82 -10 -75

rect 7 -99 24 -25

rect 184 -33 189 -25

rect 206 -33 210 -16

rect 184 -41 210 -33

rect 134 -55 161 -46

rect 134 -72 141 -55

rect 158 -72 161 -55

rect 227 -63 244 9

rect 261 -13 296 -8

rect 395 -13 412 9

rect 261 -15 412 -13

rect 261 -32 269 -15

rect 286 -30 412 -15

rect 286 -32 296 -30

rect 261 -39 296 -32

rect 261 -40 292 -39

rect 313 -56 346 -49

rect 313 -63 321 -56

rect 134 -80 161 -72

rect 178 -73 321 -63

rect 338 -73 346 -56

rect 178 -80 346 -73

rect 178 -97 195 -80

rect 395 -97 412 -30

rect 453 -56 486 -48

rect 453 -73 461 -56

rect 478 -73 486 -56

rect 453 -80 486 -73

rect 504 -64 521 9

rect 616 -13 633 9

rect 793 -13 822 -12

rect 616 -20 822 -13

rect 616 -30 798 -20

rect 566 -57 599 -49

rect 566 -64 574 -57

rect 504 -74 574 -64

rect 591 -74 599 -57

rect 504 -81 599 -74

rect -53 -107 -19 -99

rect -53 -135 -43 -107

rect -26 -135 -19 -107

rect -53 -141 -19 -135

rect -2 -107 32 -99

rect -2 -135 6 -107

rect 23 -135 32 -107

rect -2 -141 32 -135

rect 64 -105 97 -97

rect 64 -133 72 -105

rect 89 -133 97 -105

rect 64 -141 97 -133

rect 164 -105 195 -97

rect 164 -133 172 -105

rect 189 -133 195 -105

rect 164 -141 195 -133

rect 264 -105 295 -97

rect 264 -133 271 -105

rect 288 -133 295 -105

rect 264 -141 295 -133

rect 333 -105 366 -97

rect 333 -133 343 -105

rect 360 -133 366 -105

rect 333 -141 366 -133

rect 383 -105 416 -97

rect 504 -99 521 -81

rect 616 -99 633 -30

rect 793 -37 798 -30

rect 815 -37 822 -20

rect 793 -45 822 -37

rect 685 -55 719 -49

rect 685 -56 695 -55

rect 685 -73 694 -56

rect 712 -72 719 -55

rect 711 -73 719 -72

rect 685 -80 719 -73

rect 743 -55 770 -47

rect 743 -72 748 -55

rect 765 -72 770 -55

rect 839 -63 856 9

rect 874 -13 902 -8

rect 1004 -13 1021 9

rect 874 -16 1021 -13

rect 874 -33 879 -16

rect 896 -30 1021 -16

rect 896 -33 902 -30

rect 874 -41 902 -33

rect 922 -56 955 -49

rect 922 -63 930 -56

rect 743 -80 770 -72

rect 787 -73 930 -63

rect 947 -73 955 -56

rect 787 -80 955 -73

rect 787 -97 804 -80

rect 1004 -97 1021 -30

rect 383 -133 392 -105

rect 409 -133 416 -105

rect 383 -141 416 -133

rect 444 -107 478 -99

rect 444 -135 454 -107

rect 471 -135 478 -107

rect 444 -141 478 -135

rect 495 -107 529 -99

rect 495 -135 503 -107

rect 520 -135 529 -107

rect 495 -141 529 -135

rect 556 -107 590 -99

rect 556 -135 566 -107

rect 583 -135 590 -107

rect 556 -141 590 -135

rect 607 -107 641 -99

rect 607 -135 615 -107

rect 632 -135 641 -107

rect 607 -141 641 -135

rect 673 -105 706 -97

rect 673 -133 681 -105

rect 698 -133 706 -105

rect 673 -141 706 -133

rect 773 -105 804 -97

rect 773 -133 781 -105

rect 798 -133 804 -105

rect 773 -141 804 -133

rect 873 -105 904 -97

rect 873 -133 880 -105

rect 897 -133 904 -105

rect 873 -141 904 -133

rect 942 -105 975 -97

rect 942 -133 952 -105

rect 969 -133 975 -105

rect 942 -141 975 -133

rect 992 -105 1025 -97

rect 992 -133 1001 -105

rect 1018 -133 1025 -105

rect 992 -141 1025 -133

rect -43 -168 -26 -141

rect 71 -168 88 -141

rect 270 -168 287 -141

rect 343 -168 360 -141

rect 454 -168 471 -141

rect 566 -168 583 -141

rect 680 -168 697 -141

rect 879 -168 896 -141

rect 952 -168 969 -141

rect -101 -173 1051 -168

rect -101 -191 -83 -173

rect -66 -191 -42 -173

rect -25 -191 -10 -173

rect 7 -191 28 -173

rect 45 -191 71 -173

rect 88 -191 108 -173

rect 125 -191 151 -173

rect 168 -191 194 -173

rect 211 -191 237 -173

rect 254 -191 269 -173

rect 286 -191 305 -173

rect 322 -191 343 -173

rect 360 -191 373 -173

rect 390 -191 414 -173

rect 431 -191 455 -173

rect 472 -191 487 -173

rect 504 -191 525 -173

rect 542 -191 567 -173

rect 584 -191 599 -173

rect 616 -191 637 -173

rect 654 -191 680 -173

rect 697 -191 717 -173

rect 734 -191 760 -173

rect 777 -191 803 -173

rect 820 -191 846 -173

rect 863 -191 878 -173

rect 895 -191 914 -173

rect 931 -191 952 -173

rect 969 -191 996 -173

rect 1013 -191 1051 -173

rect -101 -197 1051 -191

<< viali >>

rect -82 101 -65 119

rect -46 101 -29 119

rect 122 104 139 122

rect 343 104 360 122

rect 415 101 432 119

rect 451 101 468 119

rect 563 101 580 119

rect 731 104 748 122

rect 952 104 969 122

rect 71 16 88 45

rect 172 17 189 46

rect 274 17 291 46

rect 680 16 697 45

rect 781 17 798 46

rect 883 17 900 46

rect -38 -75 -35 -58

rect -35 -75 -21 -58

rect 141 -72 158 -55

rect 461 -73 478 -56

rect 574 -74 591 -57

rect 695 -56 712 -55

rect 695 -72 711 -56

rect 711 -72 712 -56

rect 748 -72 765 -55

rect 392 -133 409 -108

rect -83 -191 -66 -173

rect -42 -191 -25 -173

rect 71 -191 88 -173

rect 269 -191 286 -173

rect 343 -191 360 -173

rect 414 -191 431 -173

rect 455 -191 472 -173

rect 567 -191 584 -173

rect 680 -191 697 -173

rect 878 -191 895 -173

rect 952 -191 969 -173

<< metal1 >>

rect -95 122 1051 125

rect -95 119 122 122

rect -95 101 -82 119

rect -65 101 -46 119

rect -29 104 122 119

rect 139 104 343 122

rect 360 119 731 122

rect 360 104 415 119

rect -29 101 415 104

rect 432 101 451 119

rect 468 101 563 119

rect 580 104 731 119

rect 748 104 952 122

rect 969 104 1051 122

rect 580 101 1051 104

rect -95 96 1051 101

rect 63 45 97 53

rect 63 16 71 45

rect 88 38 97 45

rect 164 46 197 53

rect 164 38 172 46

rect 88 20 172 38

rect 88 16 97 20

rect 63 9 97 16

rect 164 17 172 20

rect 189 38 197 46

rect 264 46 301 53

rect 264 38 274 46

rect 189 20 274 38

rect 189 17 197 20

rect 164 9 197 17

rect 264 17 274 20

rect 291 17 301 46

rect 264 9 301 17

rect 672 45 706 53

rect 672 16 680 45

rect 697 38 706 45

rect 773 46 806 53

rect 773 38 781 46

rect 697 20 781 38

rect 697 16 706 20

rect 672 9 706 16

rect 773 17 781 20

rect 798 38 806 46

rect 873 46 910 53

rect 873 38 883 46

rect 798 20 883 38

rect 798 17 806 20

rect 773 9 806 17

rect 873 17 883 20

rect 900 17 910 46

rect 873 9 910 17

rect -42 -58 -9 -51

rect -42 -75 -38 -58

rect -21 -63 -9 -58

rect 134 -55 161 -46

rect 134 -63 141 -55

rect -21 -72 141 -63

rect 158 -59 161 -55

rect 456 -56 487 -48

rect 456 -59 461 -56

rect 158 -72 461 -59

rect -21 -73 461 -72

rect 478 -73 487 -56

rect -21 -75 161 -73

rect -42 -77 161 -75

rect -42 -84 -9 -77

rect 134 -80 161 -77

rect 456 -80 487 -73

rect 563 -52 602 -47

rect 563 -79 568 -52

rect 597 -79 602 -52

rect 563 -83 602 -79

rect 688 -55 720 -47

rect 688 -72 695 -55

rect 712 -72 720 -55

rect 688 -82 720 -72

rect 737 -51 776 -47

rect 737 -78 743 -51

rect 772 -78 776 -51

rect 387 -108 412 -99

rect 387 -133 392 -108

rect 409 -116 412 -108

rect 692 -116 708 -82

rect 737 -83 776 -78

rect 409 -131 708 -116

rect 409 -133 412 -131

rect 387 -140 412 -133

rect -101 -173 1051 -168

rect -101 -191 -83 -173

rect -66 -191 -42 -173

rect -25 -191 71 -173

rect 88 -191 269 -173

rect 286 -191 343 -173

rect 360 -191 414 -173

rect 431 -191 455 -173

rect 472 -191 567 -173

rect 584 -191 680 -173

rect 697 -191 878 -173

rect 895 -191 952 -173

rect 969 -191 1051 -173

rect -101 -197 1051 -191

<< via1 >>

rect 568 -57 597 -52

rect 568 -74 574 -57

rect 574 -74 591 -57

rect 591 -74 597 -57

rect 568 -79 597 -74

rect 743 -55 772 -51

rect 743 -72 748 -55

rect 748 -72 765 -55

rect 765 -72 772 -55

rect 743 -78 772 -72

<< metal2 >>

rect 563 -52 602 -47

rect 563 -79 568 -52

rect 597 -60 602 -52

rect 737 -51 776 -47

rect 737 -60 743 -51

rect 597 -75 743 -60

rect 597 -79 602 -75

rect 563 -83 602 -79

rect 737 -78 743 -75

rect 772 -78 776 -51

rect 737 -83 776 -78

<< labels >>

flabel locali s -95 98 -61 122 0 FreeSans 80 0 0 0 VDD

port 0 nsew

flabel locali s -96 -194 -62 -170 0 FreeSans 80 0 0 0 GND

port 1 nsew

flabel poly s 86 -53 120 -29 0 FreeSans 80 0 0 0 D

port 2 nsew

flabel poly s -29 -37 5 -13 0 FreeSans 80 0 0 0 CLK

port 3 nsew

flabel locali s 995 -81 1029 -57 0 FreeSans 80 0 0 0 Q

port 4 nsew

<< end >>
