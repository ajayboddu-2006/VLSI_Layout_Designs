* SPICE3 file created from Half_Adder.ext - technology: sky130A
.include pshort.lib
.include nshort.lib
.option scale=0.01u

//.subckt Half_Adder VDD GND A B SUM COUT
M1000 COUT a_494_9# VDD VDD pshort_model.0 ad=1620 pd=162 as=1490 ps=156 w=45 l=15
M1001 a_494_9# B a_494_n141# GND nshort_model.0 ad=1540 pd=158 as=770 ps=79u w=44 l=15
M1002 a_n117_n141# A VDD VDD pshort_model.0 ad=1670 pd=164 as=1620 ps=162 w=45 l=15
M1003 a_n3_n147# B VDD VDD pshort_model.0 ad=1540 pd=158 as=1540 ps=158 w=44 l=15
M1004 GND A a_213_n146# GND nshort_model.0 ad=1410 pd=152 as=770 ps=79u w=44 l=15
M1005 a_163_n146# a_n3_n147# a_63_9# VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1006 a_63_9# B VDD VDD pshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1007 a_163_n146# B a_113_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1008 VDD a_n117_n141# a_63_9# VDD pshort_model.0 ad=770 pd=79u as=1540 ps=158 w=44 l=15
M1009 a_494_9# A VDD VDD pshort_model.0 ad=787 pd=80u as=1580 ps=160 w=45 l=15
M1010 COUT a_494_9# GND GND nshort_model.0 ad=1500 pd=156 as=1450 ps=154 w=44 l=15
M1011 a_63_9# A a_163_n146# VDD pshort_model.0 ad=1670 pd=164 as=770 ps=79u w=44 l=15
M1012 a_n117_n141# A GND GND nshort_model.0 ad=1510 pd=156 as=1510 ps=156 w=42 l=15
M1013 a_113_n146# a_n117_n141# GND GND nshort_model.0 ad=770 pd=79u as=1500 ps=156 w=44 l=15
M1014 a_494_n141# A GND GND nshort_model.0 ad=770 pd=79u as=1450 ps=154 w=44 l=15
M1015 a_n3_n147# B GND GND nshort_model.0 ad=1580 pd=160 as=1580 ps=160 w=45 l=15
M1016 VDD B a_494_9# VDD pshort_model.0 ad=1580 pd=79u as=787 ps=80u w=45 l=15
M1017 SUM a_163_n146# GND GND nshort_model.0 ad=1500 pd=156 as=1500 ps=156 w=44 l=15
M1018 a_213_n146# a_n3_n147# a_163_n146# GND nshort_model.0 ad=770 pd=79u as=770 ps=79u w=44 l=15
M1019 SUM a_163_n146# VDD VDD pshort_model.0 ad=1580 pd=160 as=1530 ps=158 w=45 l=15

VDD VDD 0 5V
VSS VSS 0 0V
Va A VSS PULSE(0 5V 0 0.1ns 0.1ns 5ns 10ns)
Vb B VSS PULSE(0 5V 0 0.1ns 0.1ns 4ns 8ns)

C0 VDD B 0.0473f
C1 VDD a_n3_n147# 0.188f
C2 A B 0.127f
C3 a_n3_n147# A 0.096f
C4 VDD A 0.0432f
C5 a_494_9# SUM 0.0393f
C6 a_163_n146# a_113_n146# 0.00374f
C7 a_163_n146# a_213_n146# 0.00731f
C8 a_n3_n147# a_113_n146# 0.00282f
C9 a_494_9# B 0.0812f
C10 VDD a_494_n141# 1.69e-19
C11 VDD a_494_9# 0.263f
C12 A a_494_9# 0.0187f
C13 SUM a_63_9# 0.00219f
C14 COUT B 7.94e-19
C15 VDD COUT 0.126f
C16 a_163_n146# a_63_9# 0.228f
C17 a_n117_n141# a_63_9# 0.0253f
C18 B a_63_9# 0.0137f
C19 a_n3_n147# a_63_9# 0.163f
C20 a_163_n146# SUM 0.0574f
C21 VDD a_63_9# 0.551f
C22 a_494_9# a_494_n141# 0.00699f
C23 A a_63_9# 0.0136f
C24 a_n117_n141# a_163_n146# 0.0157f
C25 SUM B 2.46e-19
C26 a_n3_n147# SUM 1.16e-19
C27 a_494_9# COUT 0.0646f
C28 VDD SUM 0.183f
C29 a_163_n146# B 0.0107f
C30 A SUM 0.00716f
C31 a_n3_n147# a_163_n146# 0.171f
C32 VDD a_163_n146# 0.0681f
C33 a_n117_n141# B 0.158f
C34 a_n3_n147# a_n117_n141# 0.229f
C35 a_163_n146# A 0.105f
C36 a_63_9# a_113_n146# 0.00134f
C37 VDD a_n117_n141# 0.238f
C38 a_213_n146# a_63_9# 0.00134f
C39 a_n117_n141# A 0.025f
C40 a_494_9# a_63_9# 1.36e-19
C41 a_n3_n147# B 0.152f
C42 COUT GND 0.272f
C43 SUM GND 0.253f
C44 B GND 0.511f
C45 A GND 0.578f
C46 VDD GND 3.23f
C47 a_494_n141# GND 0.0088f **FLOATING
C48 a_213_n146# GND 0.00892f **FLOATING
C49 a_113_n146# GND 0.00892f **FLOATING
C50 a_63_9# GND 0.135f **FLOATING
C51 a_494_9# GND 0.548f **FLOATING
C52 a_163_n146# GND 0.578f **FLOATING
C53 a_n3_n147# GND 0.481f **FLOATING
C54 a_n117_n141# GND 0.746f **FLOATING
//.ends
.tran 1n 20n
.control
run
.endc
.end
