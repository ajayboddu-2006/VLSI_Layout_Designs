magic
tech sky130A
timestamp 1737026182
<< nwell >>
rect -86 148 115 290
<< nmos >>
rect -27 34 -12 82
rect 24 34 39 82
<< pmos >>
rect -27 166 -12 211
rect 24 166 39 211
<< ndiff >>
rect -64 74 -27 82
rect -64 42 -55 74
rect -34 42 -27 74
rect -64 34 -27 42
rect -12 34 24 82
rect 39 74 78 82
rect 39 42 49 74
rect 70 42 78 74
rect 39 34 78 42
<< pdiff >>
rect -62 204 -27 211
rect -62 173 -54 204
rect -37 173 -27 204
rect -62 166 -27 173
rect -12 204 24 211
rect -12 173 -2 204
rect 15 173 24 204
rect -12 166 24 173
rect 39 204 72 211
rect 39 173 48 204
rect 65 173 72 204
rect 39 166 72 173
<< ndiffc >>
rect -55 42 -34 74
rect 49 42 70 74
<< pdiffc >>
rect -54 173 -37 204
rect -2 173 15 204
rect 48 173 65 204
<< psubdiff >>
rect -94 -27 107 -24
rect -94 -44 -80 -27
rect -63 -28 78 -27
rect -63 -44 -25 -28
rect -94 -45 -25 -44
rect -8 -45 9 -28
rect 26 -45 44 -28
rect 61 -44 78 -28
rect 95 -44 107 -27
rect 61 -45 107 -44
rect -94 -49 107 -45
<< nsubdiff >>
rect -68 269 90 272
rect -68 268 36 269
rect -68 251 -34 268
rect -17 251 0 268
rect 17 252 36 268
rect 53 252 90 269
rect 17 251 90 252
rect -68 247 90 251
<< psubdiffcont >>
rect -80 -44 -63 -27
rect -25 -45 -8 -28
rect 9 -45 26 -28
rect 44 -45 61 -28
rect 78 -44 95 -27
<< nsubdiffcont >>
rect -34 251 -17 268
rect 0 251 17 268
rect 36 252 53 269
<< poly >>
rect -27 211 -12 233
rect 24 211 39 233
rect -89 137 -58 145
rect -89 120 -80 137
rect -63 135 -58 137
rect -27 135 -12 166
rect -63 120 -12 135
rect -89 112 -58 120
rect -27 82 -12 120
rect 24 143 39 166
rect 75 143 114 149
rect 24 139 114 143
rect 24 124 87 139
rect 24 82 39 124
rect 75 122 87 124
rect 104 122 114 139
rect 75 112 114 122
rect -27 -8 -12 34
rect 24 -8 39 34
<< polycont >>
rect -80 120 -63 137
rect 87 122 104 139
<< locali >>
rect -86 269 114 272
rect -86 252 -63 269
rect -46 268 36 269
rect -46 252 -34 268
rect -86 251 -34 252
rect -17 251 0 268
rect 17 252 36 268
rect 53 252 55 269
rect 72 252 114 269
rect 17 251 114 252
rect -86 247 114 251
rect -62 211 -45 247
rect 55 211 72 247
rect -62 204 -29 211
rect -62 173 -54 204
rect -37 173 -29 204
rect -62 166 -29 173
rect -10 204 23 211
rect -10 173 -2 204
rect 15 173 23 204
rect -10 166 23 173
rect 40 204 73 211
rect 40 173 48 204
rect 65 173 73 204
rect 40 166 73 173
rect -89 137 -58 145
rect -97 120 -80 137
rect -63 120 -58 137
rect -89 112 -58 120
rect -2 113 15 166
rect 75 141 114 149
rect 75 139 120 141
rect 75 122 87 139
rect 104 122 120 139
rect 75 121 120 122
rect -2 96 58 113
rect 75 112 114 121
rect 41 82 58 96
rect -64 74 -28 82
rect -64 42 -55 74
rect -34 42 -28 74
rect -64 34 -28 42
rect 41 74 78 82
rect 41 42 49 74
rect 70 42 78 74
rect 41 34 78 42
rect -57 -24 -39 34
rect -94 -27 107 -24
rect -94 -44 -80 -27
rect -63 -28 78 -27
rect -63 -44 -56 -28
rect -94 -45 -56 -44
rect -39 -45 -25 -28
rect -8 -45 9 -28
rect 26 -45 44 -28
rect 61 -44 78 -28
rect 95 -44 107 -27
rect 61 -45 107 -44
rect -94 -49 107 -45
<< viali >>
rect -63 252 -46 269
rect 55 252 72 269
rect -56 -45 -39 -28
<< metal1 >>
rect -86 269 114 272
rect -86 252 -63 269
rect -46 252 55 269
rect 72 252 114 269
rect -86 247 114 252
rect -94 -28 107 -24
rect -94 -45 -56 -28
rect -39 -45 107 -28
rect -94 -49 107 -45
<< labels >>
flabel space -89 248 -62 269 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel metal1 -93 -47 -66 -26 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel locali -88 115 -61 136 0 FreeSans 80 0 0 0 IN1
port 2 nsew
flabel locali 81 123 108 144 0 FreeSans 80 0 0 0 IN2
port 3 nsew
flabel space 33 96 60 117 0 FreeSans 80 0 0 0 OUT
port 4 nsew
<< end >>
