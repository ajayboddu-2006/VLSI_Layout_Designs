magic

tech sky130A

timestamp 1737430450

<< nwell >>

rect -191 -15 708 143

<< nmos >>

rect -132 -141 -117 -99

rect -18 -147 -3 -102

rect 98 -146 113 -102

rect 148 -146 163 -102

rect 198 -146 213 -102

rect 248 -146 263 -102

rect 367 -141 382 -97

rect 479 -141 494 -97

rect 529 -141 544 -97

rect 639 -141 654 -97

<< pmos >>

rect -132 9 -117 54

rect -18 9 -3 53

rect 98 9 113 53

rect 148 9 163 53

rect 198 9 213 53

rect 248 9 263 53

rect 367 9 382 54

rect 479 9 494 54

rect 529 9 544 54

rect 639 9 654 54

<< ndiff >>

rect -168 -105 -132 -99

rect -168 -133 -159 -105

rect -142 -133 -132 -105

rect -168 -141 -132 -133

rect -117 -105 -81 -99

rect -117 -133 -106 -105

rect -89 -133 -81 -105

rect -117 -141 -81 -133

rect -53 -110 -18 -102

rect -53 -138 -43 -110

rect -26 -138 -18 -110

rect -53 -147 -18 -138

rect -3 -110 32 -102

rect -3 -138 6 -110

rect 23 -138 32 -110

rect -3 -147 32 -138

rect 64 -109 98 -102

rect 64 -137 72 -109

rect 89 -137 98 -109

rect 64 -146 98 -137

rect 113 -146 148 -102

rect 163 -110 198 -102

rect 163 -138 172 -110

rect 189 -138 198 -110

rect 163 -146 198 -138

rect 213 -146 248 -102

rect 263 -110 295 -102

rect 263 -138 271 -110

rect 288 -138 295 -110

rect 263 -146 295 -138

rect 333 -105 367 -97

rect 333 -133 343 -105

rect 360 -133 367 -105

rect 333 -141 367 -133

rect 382 -105 416 -97

rect 382 -133 392 -105

rect 409 -133 416 -105

rect 382 -141 416 -133

rect 446 -105 479 -97

rect 446 -133 454 -105

rect 471 -133 479 -105

rect 446 -141 479 -133

rect 494 -141 529 -97

rect 544 -105 579 -97

rect 544 -133 553 -105

rect 570 -133 579 -105

rect 544 -141 579 -133

rect 606 -105 639 -97

rect 606 -133 614 -105

rect 631 -133 639 -105

rect 606 -141 639 -133

rect 654 -105 688 -97

rect 654 -133 664 -105

rect 681 -133 688 -105

rect 654 -141 688 -133

<< pdiff >>

rect -168 46 -132 54

rect -168 17 -160 46

rect -142 17 -132 46

rect -168 9 -132 17

rect -117 45 -80 54

rect -117 16 -107 45

rect -89 16 -80 45

rect -117 9 -80 16

rect -53 46 -18 53

rect -53 17 -45 46

rect -27 17 -18 46

rect -53 9 -18 17

rect -3 46 32 53

rect -3 17 6 46

rect 24 17 32 46

rect -3 9 32 17

rect 63 45 98 53

rect 63 16 71 45

rect 89 16 98 45

rect 63 9 98 16

rect 113 45 148 53

rect 113 16 122 45

rect 139 16 148 45

rect 113 9 148 16

rect 163 46 198 53

rect 163 17 172 46

rect 189 17 198 46

rect 163 9 198 17

rect 213 46 248 53

rect 213 17 222 46

rect 239 17 248 46

rect 213 9 248 17

rect 263 46 301 53

rect 263 17 274 46

rect 291 17 301 46

rect 263 9 301 17

rect 333 46 367 54

rect 333 17 342 46

rect 359 17 367 46

rect 333 9 367 17

rect 382 45 417 54

rect 382 16 392 45

rect 409 16 417 45

rect 382 9 417 16

rect 444 46 479 54

rect 444 17 451 46

rect 468 17 479 46

rect 444 9 479 17

rect 494 47 529 54

rect 494 18 503 47

rect 520 18 529 47

rect 494 9 529 18

rect 544 47 579 54

rect 544 18 554 47

rect 571 18 579 47

rect 544 9 579 18

rect 606 46 639 54

rect 606 17 614 46

rect 631 17 639 46

rect 606 9 639 17

rect 654 47 690 54

rect 654 18 665 47

rect 682 18 690 47

rect 654 9 690 18

<< ndiffc >>

rect -159 -133 -142 -105

rect -106 -133 -89 -105

rect -43 -138 -26 -110

rect 6 -138 23 -110

rect 72 -137 89 -109

rect 172 -138 189 -110

rect 271 -138 288 -110

rect 343 -133 360 -105

rect 392 -133 409 -105

rect 454 -133 471 -105

rect 553 -133 570 -105

rect 614 -133 631 -105

rect 664 -133 681 -105

<< pdiffc >>

rect -160 17 -142 46

rect -107 16 -89 45

rect -45 17 -27 46

rect 6 17 24 46

rect 71 16 89 45

rect 122 16 139 45

rect 172 17 189 46

rect 222 17 239 46

rect 274 17 291 46

rect 342 17 359 46

rect 392 16 409 45

rect 451 17 468 46

rect 503 18 520 47

rect 554 18 571 47

rect 614 17 631 46

rect 665 18 682 47

<< psubdiff >>

rect -189 -190 698 -186

rect -189 -208 -122 -190

rect -105 -191 422 -190

rect -105 -208 -10 -191

rect -189 -209 -10 -208

rect 7 -209 28 -191

rect 45 -209 108 -191

rect 125 -209 151 -191

rect 168 -209 194 -191

rect 211 -209 237 -191

rect 254 -209 305 -191

rect 322 -209 387 -191

rect 404 -208 422 -191

rect 439 -191 698 -190

rect 439 -208 490 -191

rect 404 -209 490 -208

rect 507 -209 532 -191

rect 549 -209 574 -191

rect 591 -209 659 -191

rect 676 -209 698 -191

rect -189 -215 698 -209

<< nsubdiff >>

rect -173 122 685 125

rect -173 121 379 122

rect -173 103 -122 121

rect -105 119 24 121

rect -105 103 -12 119

rect -173 101 -12 103

rect 5 103 24 119

rect 41 120 94 121

rect 41 103 60 120

rect 5 102 60 103

rect 77 103 94 120

rect 111 103 162 121

rect 179 120 313 121

rect 179 103 200 120

rect 77 102 200 103

rect 217 119 276 120

rect 217 102 240 119

rect 5 101 240 102

rect 257 102 276 119

rect 293 103 313 120

rect 330 104 379 121

rect 396 104 417 122

rect 434 121 685 122

rect 434 120 586 121

rect 434 104 491 120

rect 330 103 491 104

rect 293 102 491 103

rect 508 102 527 120

rect 544 103 586 120

rect 603 103 642 121

rect 659 103 685 121

rect 544 102 685 103

rect 257 101 685 102

rect -173 96 685 101

<< psubdiffcont >>

rect -122 -208 -105 -190

rect -10 -209 7 -191

rect 28 -209 45 -191

rect 108 -209 125 -191

rect 151 -209 168 -191

rect 194 -209 211 -191

rect 237 -209 254 -191

rect 305 -209 322 -191

rect 387 -209 404 -191

rect 422 -208 439 -190

rect 490 -209 507 -191

rect 532 -209 549 -191

rect 574 -209 591 -191

rect 659 -209 676 -191

<< nsubdiffcont >>

rect -122 103 -105 121

rect -12 101 5 119

rect 24 103 41 121

rect 60 102 77 120

rect 94 103 111 121

rect 162 103 179 121

rect 200 102 217 120

rect 240 101 257 119

rect 276 102 293 120

rect 313 103 330 121

rect 379 104 396 122

rect 417 104 434 122

rect 491 102 508 120

rect 527 102 544 120

rect 586 103 603 121

rect 642 103 659 121

<< poly >>

rect -132 54 -117 75

rect -18 53 -3 75

rect 98 53 113 75

rect 148 53 163 75

rect 198 53 213 75

rect 248 53 263 75

rect 367 54 382 75

rect 479 54 494 79

rect 529 54 544 79

rect 639 54 654 79

rect -132 -99 -117 9

rect -18 -102 -3 9

rect 44 -61 77 -54

rect 98 -61 113 9

rect 44 -78 52 -61

rect 69 -76 113 -61

rect 69 -78 77 -76

rect 44 -85 77 -78

rect 98 -102 113 -76

rect 148 -102 163 9

rect 198 -12 213 9

rect 184 -20 213 -12

rect 184 -37 189 -20

rect 206 -37 213 -20

rect 184 -45 213 -37

rect 198 -102 213 -45

rect 248 -102 263 9

rect 313 -56 346 -49

rect 313 -73 321 -56

rect 338 -63 346 -56

rect 367 -63 382 9

rect 338 -73 382 -63

rect 313 -80 382 -73

rect 367 -97 382 -80

rect 479 -97 494 9

rect 529 -97 544 9

rect 585 -55 618 -49

rect 585 -72 593 -55

rect 610 -63 618 -55

rect 639 -63 654 9

rect 610 -72 654 -63

rect 585 -80 654 -72

rect 639 -97 654 -80

rect -132 -158 -117 -141

rect -18 -160 -3 -147

rect 98 -159 113 -146

rect 148 -159 163 -146

rect 198 -159 213 -146

rect 248 -159 263 -146

rect 367 -154 382 -141

rect 479 -154 494 -141

rect 529 -154 544 -141

rect 639 -154 654 -141

<< polycont >>

rect 52 -78 69 -61

rect 189 -37 206 -20

rect 321 -73 338 -56

rect 593 -72 610 -55

<< locali >>

rect -191 122 703 125

rect -191 121 122 122

rect -191 103 -161 121

rect -144 103 -122 121

rect -105 119 24 121

rect -105 103 -82 119

rect -191 101 -82 103

rect -65 101 -46 119

rect -29 101 -12 119

rect 5 103 24 119

rect 41 120 94 121

rect 41 103 60 120

rect 5 102 60 103

rect 77 103 94 120

rect 111 104 122 121

rect 139 121 343 122

rect 139 104 162 121

rect 111 103 162 104

rect 179 120 313 121

rect 179 103 200 120

rect 77 102 200 103

rect 217 119 276 120

rect 217 102 240 119

rect 5 101 240 102

rect 257 102 276 119

rect 293 103 313 120

rect 330 104 343 121

rect 360 104 379 122

rect 396 104 417 122

rect 434 121 703 122

rect 434 120 586 121

rect 434 104 451 120

rect 330 103 451 104

rect 293 102 451 103

rect 468 102 491 120

rect 508 102 527 120

rect 544 102 552 120

rect 569 103 586 120

rect 603 120 642 121

rect 603 103 613 120

rect 569 102 613 103

rect 630 103 642 120

rect 659 103 703 121

rect 630 102 703 103

rect 257 101 703 102

rect -191 96 703 101

rect -162 54 -143 96

rect -168 46 -134 54

rect -168 17 -160 46

rect -142 17 -134 46

rect -168 9 -134 17

rect -115 45 -80 54

rect -43 53 -26 96

rect 123 53 140 96

rect 344 54 361 96

rect 451 54 468 96

rect 554 54 571 96

rect 614 54 631 96

rect -115 16 -107 45

rect -89 16 -80 45

rect -115 9 -80 16

rect -53 46 -19 53

rect -53 17 -45 46

rect -27 17 -19 46

rect -53 9 -19 17

rect -2 46 32 53

rect -2 17 6 46

rect 24 17 32 46

rect -2 9 32 17

rect 63 45 97 53

rect 63 16 71 45

rect 89 16 97 45

rect 63 9 97 16

rect 114 45 147 53

rect 114 16 122 45

rect 139 16 147 45

rect 114 9 147 16

rect 164 46 197 53

rect 164 17 172 46

rect 189 17 197 46

rect 164 9 197 17

rect 214 46 247 53

rect 214 17 222 46

rect 239 17 247 46

rect 214 9 247 17

rect 264 46 301 53

rect 264 17 274 46

rect 291 17 301 46

rect 264 9 301 17

rect 333 46 366 54

rect 333 17 342 46

rect 359 17 366 46

rect 333 9 366 17

rect 383 45 417 54

rect 383 16 392 45

rect 409 16 417 45

rect 383 9 417 16

rect 444 46 478 54

rect 444 17 451 46

rect 468 17 478 46

rect 444 9 478 17

rect 495 47 528 54

rect 495 18 503 47

rect 520 18 528 47

rect 495 9 528 18

rect 545 47 579 54

rect 545 18 554 47

rect 571 18 579 47

rect 545 9 579 18

rect 606 46 638 54

rect 606 17 614 46

rect 631 17 638 46

rect 606 9 638 17

rect 655 47 690 54

rect 655 18 665 47

rect 682 18 690 47

rect 655 9 690 18

rect -107 -63 -89 9

rect 7 -20 24 9

rect 184 -20 213 -12

rect 7 -37 189 -20

rect 206 -37 213 -20

rect -62 -63 -32 -57

rect -107 -80 -55 -63

rect -38 -80 -32 -63

rect -107 -99 -89 -80

rect -62 -85 -32 -80

rect -168 -105 -134 -99

rect -168 -133 -159 -105

rect -142 -133 -134 -105

rect -168 -141 -134 -133

rect -115 -105 -81 -99

rect 7 -102 24 -37

rect 184 -45 213 -37

rect 44 -61 77 -54

rect 44 -78 52 -61

rect 69 -78 77 -61

rect 230 -63 247 9

rect 395 -40 412 9

rect 313 -56 346 -49

rect 313 -63 321 -56

rect 44 -85 77 -78

rect 171 -73 321 -63

rect 338 -73 346 -56

rect 171 -80 346 -73

rect 395 -57 439 -40

rect 171 -102 188 -80

rect 395 -97 412 -57

rect 502 -63 519 9

rect 665 -43 682 9

rect 585 -55 618 -49

rect 585 -63 593 -55

rect 502 -72 593 -63

rect 610 -72 618 -55

rect 502 -80 618 -72

rect 665 -60 706 -43

rect 553 -97 570 -80

rect 665 -97 682 -60

rect -115 -133 -106 -105

rect -89 -133 -81 -105

rect -115 -141 -81 -133

rect -53 -110 -19 -102

rect -53 -138 -43 -110

rect -26 -138 -19 -110

rect -159 -186 -142 -141

rect -53 -147 -19 -138

rect -2 -110 32 -102

rect -2 -138 6 -110

rect 23 -138 32 -110

rect -2 -147 32 -138

rect 64 -109 97 -102

rect 64 -137 72 -109

rect 89 -137 97 -109

rect 64 -146 97 -137

rect 164 -110 195 -102

rect 164 -138 172 -110

rect 189 -138 195 -110

rect 164 -146 195 -138

rect 264 -110 295 -102

rect 264 -138 271 -110

rect 288 -138 295 -110

rect 264 -146 295 -138

rect 333 -105 366 -97

rect 333 -133 343 -105

rect 360 -133 366 -105

rect 333 -141 366 -133

rect 383 -105 416 -97

rect 383 -133 392 -105

rect 409 -133 416 -105

rect 383 -141 416 -133

rect 446 -105 478 -97

rect 446 -133 454 -105

rect 471 -133 478 -105

rect 446 -141 478 -133

rect 545 -105 579 -97

rect 545 -133 553 -105

rect 570 -133 579 -105

rect 545 -141 579 -133

rect 606 -105 638 -97

rect 606 -133 614 -105

rect 631 -133 638 -105

rect 606 -141 638 -133

rect 656 -105 688 -97

rect 656 -133 664 -105

rect 681 -133 688 -105

rect 656 -141 688 -133

rect -43 -186 -26 -147

rect 71 -186 88 -146

rect 270 -186 287 -146

rect 343 -186 360 -141

rect 454 -186 471 -141

rect 614 -186 631 -141

rect -189 -190 698 -186

rect -189 -191 -122 -190

rect -189 -209 -160 -191

rect -143 -208 -122 -191

rect -105 -191 422 -190

rect -105 -208 -83 -191

rect -143 -209 -83 -208

rect -66 -209 -42 -191

rect -25 -209 -10 -191

rect 7 -209 28 -191

rect 45 -209 71 -191

rect 88 -209 108 -191

rect 125 -209 151 -191

rect 168 -209 194 -191

rect 211 -209 237 -191

rect 254 -209 269 -191

rect 286 -209 305 -191

rect 322 -209 343 -191

rect 360 -209 387 -191

rect 404 -208 422 -191

rect 439 -191 614 -190

rect 439 -208 454 -191

rect 404 -209 454 -208

rect 471 -209 490 -191

rect 507 -209 532 -191

rect 549 -209 574 -191

rect 591 -208 614 -191

rect 631 -191 698 -190

rect 631 -208 659 -191

rect 591 -209 659 -208

rect 676 -209 698 -191

rect -189 -215 698 -209

<< viali >>

rect -161 103 -144 121

rect -82 101 -65 119

rect -46 101 -29 119

rect 122 104 139 122

rect 343 104 360 122

rect 451 102 468 120

rect 552 102 569 120

rect 613 102 630 120

rect 71 16 88 45

rect 172 17 189 46

rect 274 17 291 46

rect -55 -80 -38 -63

rect 52 -78 69 -61

rect -160 -209 -143 -191

rect -83 -209 -66 -191

rect -42 -209 -25 -191

rect 71 -209 88 -191

rect 269 -209 286 -191

rect 343 -209 360 -191

rect 454 -209 471 -191

rect 614 -208 631 -190

<< metal1 >>

rect -191 122 703 125

rect -191 121 122 122

rect -191 103 -161 121

rect -144 119 122 121

rect -144 103 -82 119

rect -191 101 -82 103

rect -65 101 -46 119

rect -29 104 122 119

rect 139 104 343 122

rect 360 120 703 122

rect 360 104 451 120

rect -29 102 451 104

rect 468 102 552 120

rect 569 102 613 120

rect 630 102 703 120

rect -29 101 703 102

rect -191 96 703 101

rect 63 45 97 53

rect 63 16 71 45

rect 88 38 97 45

rect 164 46 197 53

rect 164 38 172 46

rect 88 20 172 38

rect 88 16 97 20

rect 63 9 97 16

rect 164 17 172 20

rect 189 38 197 46

rect 264 46 301 53

rect 264 38 274 46

rect 189 20 274 38

rect 189 17 197 20

rect 164 9 197 17

rect 264 17 274 20

rect 291 17 301 46

rect 264 9 301 17

rect -62 -63 -32 -57

rect 44 -61 77 -54

rect 44 -63 52 -61

rect -62 -80 -55 -63

rect -38 -78 52 -63

rect 69 -78 77 -61

rect -38 -80 -32 -78

rect -62 -85 -32 -80

rect 44 -85 77 -78

rect -189 -190 698 -186

rect -189 -191 614 -190

rect -189 -209 -160 -191

rect -143 -209 -83 -191

rect -66 -209 -42 -191

rect -25 -209 71 -191

rect 88 -209 269 -191

rect 286 -209 343 -191

rect 360 -209 454 -191

rect 471 -208 614 -191

rect 631 -208 698 -190

rect 471 -209 698 -208

rect -189 -215 698 -209

<< labels >>

flabel metal1 s -189 100 -165 120 0 FreeSans 80 0 0 0 VDD

port 0 nsew

flabel metal1 s -187 -211 -163 -191 0 FreeSans 80 0 0 0 GND

port 1 nsew

flabel poly s -138 -163 -114 -143 0 FreeSans 80 0 0 0 A

port 2 nsew

flabel poly s 243 -167 267 -147 0 FreeSans 80 0 0 0 A

flabel poly s -21 -167 3 -147 0 FreeSans 80 0 0 0 B

port 3 nsew

flabel poly s 144 -167 168 -147 0 FreeSans 80 0 0 0 B

flabel poly s 475 -155 498 -142 0 FreeSans 80 0 0 0 A

flabel poly s 527 -156 550 -143 0 FreeSans 80 0 0 0 B

flabel locali s 416 -57 439 -44 0 FreeSans 80 0 0 0 SUM

port 4 nsew

flabel locali s 666 -59 689 -46 0 FreeSans 80 0 0 0 COUT

port 5 nsew

<< end >>
