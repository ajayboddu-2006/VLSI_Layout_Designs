magic
tech sky130A
timestamp 1737465221
<< nwell >>
rect -191 -15 1893 143
<< nmos >>
rect -132 -141 -117 -99
rect -18 -147 -3 -102
rect 98 -146 113 -102
rect 148 -146 163 -102
rect 198 -146 213 -102
rect 248 -146 263 -102
rect 367 -141 382 -97
rect 479 -141 494 -97
rect 529 -141 544 -97
rect 639 -141 654 -97
rect 754 -141 769 -99
rect 868 -147 883 -102
rect 984 -146 999 -102
rect 1034 -146 1049 -102
rect 1084 -146 1099 -102
rect 1134 -146 1149 -102
rect 1253 -141 1268 -97
rect 1365 -141 1380 -97
rect 1415 -141 1430 -97
rect 1525 -141 1540 -97
rect 1639 -141 1654 -97
rect 1691 -141 1706 -97
rect 1815 -141 1830 -99
<< pmos >>
rect -132 9 -117 54
rect -18 9 -3 53
rect 98 9 113 53
rect 148 9 163 53
rect 198 9 213 53
rect 248 9 263 53
rect 367 9 382 54
rect 479 9 494 54
rect 529 9 544 54
rect 639 9 654 54
rect 754 9 769 54
rect 868 9 883 53
rect 984 9 999 53
rect 1034 9 1049 53
rect 1084 9 1099 53
rect 1134 9 1149 53
rect 1253 9 1268 54
rect 1365 9 1380 54
rect 1415 9 1430 54
rect 1525 9 1540 54
rect 1639 9 1654 54
rect 1691 9 1706 54
rect 1815 9 1830 54
<< ndiff >>
rect -168 -105 -132 -99
rect -168 -133 -159 -105
rect -142 -133 -132 -105
rect -168 -141 -132 -133
rect -117 -105 -81 -99
rect -117 -133 -106 -105
rect -89 -133 -81 -105
rect -117 -141 -81 -133
rect -53 -110 -18 -102
rect -53 -138 -43 -110
rect -26 -138 -18 -110
rect -53 -147 -18 -138
rect -3 -110 32 -102
rect -3 -138 6 -110
rect 23 -138 32 -110
rect -3 -147 32 -138
rect 64 -109 98 -102
rect 64 -137 72 -109
rect 89 -137 98 -109
rect 64 -146 98 -137
rect 113 -146 148 -102
rect 163 -110 198 -102
rect 163 -138 172 -110
rect 189 -138 198 -110
rect 163 -146 198 -138
rect 213 -146 248 -102
rect 263 -110 295 -102
rect 263 -138 271 -110
rect 288 -138 295 -110
rect 263 -146 295 -138
rect 333 -105 367 -97
rect 333 -133 343 -105
rect 360 -133 367 -105
rect 333 -141 367 -133
rect 382 -105 416 -97
rect 382 -133 392 -105
rect 409 -133 416 -105
rect 382 -141 416 -133
rect 446 -105 479 -97
rect 446 -133 454 -105
rect 471 -133 479 -105
rect 446 -141 479 -133
rect 494 -141 529 -97
rect 544 -105 579 -97
rect 544 -133 553 -105
rect 570 -133 579 -105
rect 544 -141 579 -133
rect 606 -105 639 -97
rect 606 -133 614 -105
rect 631 -133 639 -105
rect 606 -141 639 -133
rect 654 -105 688 -97
rect 654 -133 664 -105
rect 681 -133 688 -105
rect 654 -141 688 -133
rect 718 -105 754 -99
rect 718 -133 727 -105
rect 744 -133 754 -105
rect 718 -141 754 -133
rect 769 -105 805 -99
rect 769 -133 780 -105
rect 797 -133 805 -105
rect 769 -141 805 -133
rect 833 -110 868 -102
rect 833 -138 843 -110
rect 860 -138 868 -110
rect 833 -147 868 -138
rect 883 -110 918 -102
rect 883 -138 892 -110
rect 909 -138 918 -110
rect 883 -147 918 -138
rect 950 -109 984 -102
rect 950 -137 958 -109
rect 975 -137 984 -109
rect 950 -146 984 -137
rect 999 -146 1034 -102
rect 1049 -110 1084 -102
rect 1049 -138 1058 -110
rect 1075 -138 1084 -110
rect 1049 -146 1084 -138
rect 1099 -146 1134 -102
rect 1149 -110 1181 -102
rect 1149 -138 1157 -110
rect 1174 -138 1181 -110
rect 1149 -146 1181 -138
rect 1219 -105 1253 -97
rect 1219 -133 1229 -105
rect 1246 -133 1253 -105
rect 1219 -141 1253 -133
rect 1268 -105 1302 -97
rect 1268 -133 1278 -105
rect 1295 -133 1302 -105
rect 1268 -141 1302 -133
rect 1332 -105 1365 -97
rect 1332 -133 1340 -105
rect 1357 -133 1365 -105
rect 1332 -141 1365 -133
rect 1380 -141 1415 -97
rect 1430 -105 1465 -97
rect 1430 -133 1439 -105
rect 1456 -133 1465 -105
rect 1430 -141 1465 -133
rect 1492 -105 1525 -97
rect 1492 -133 1500 -105
rect 1517 -133 1525 -105
rect 1492 -141 1525 -133
rect 1540 -105 1574 -97
rect 1540 -133 1550 -105
rect 1567 -133 1574 -105
rect 1540 -141 1574 -133
rect 1605 -105 1639 -97
rect 1605 -133 1614 -105
rect 1631 -133 1639 -105
rect 1605 -141 1639 -133
rect 1654 -105 1691 -97
rect 1654 -133 1664 -105
rect 1681 -133 1691 -105
rect 1654 -141 1691 -133
rect 1706 -105 1740 -97
rect 1706 -133 1718 -105
rect 1735 -133 1740 -105
rect 1706 -141 1740 -133
rect 1779 -105 1815 -99
rect 1779 -133 1788 -105
rect 1805 -133 1815 -105
rect 1779 -141 1815 -133
rect 1830 -105 1866 -99
rect 1830 -133 1841 -105
rect 1858 -133 1866 -105
rect 1830 -141 1866 -133
<< pdiff >>
rect -168 46 -132 54
rect -168 17 -160 46
rect -142 17 -132 46
rect -168 9 -132 17
rect -117 45 -80 54
rect -117 16 -107 45
rect -89 16 -80 45
rect -117 9 -80 16
rect -53 46 -18 53
rect -53 17 -45 46
rect -27 17 -18 46
rect -53 9 -18 17
rect -3 46 32 53
rect -3 17 6 46
rect 24 17 32 46
rect -3 9 32 17
rect 63 45 98 53
rect 63 16 71 45
rect 89 16 98 45
rect 63 9 98 16
rect 113 45 148 53
rect 113 16 122 45
rect 139 16 148 45
rect 113 9 148 16
rect 163 46 198 53
rect 163 17 172 46
rect 189 17 198 46
rect 163 9 198 17
rect 213 46 248 53
rect 213 17 222 46
rect 239 17 248 46
rect 213 9 248 17
rect 263 46 301 53
rect 263 17 274 46
rect 291 17 301 46
rect 263 9 301 17
rect 333 46 367 54
rect 333 17 342 46
rect 359 17 367 46
rect 333 9 367 17
rect 382 45 417 54
rect 382 16 392 45
rect 409 16 417 45
rect 382 9 417 16
rect 444 46 479 54
rect 444 17 451 46
rect 468 17 479 46
rect 444 9 479 17
rect 494 47 529 54
rect 494 18 503 47
rect 520 18 529 47
rect 494 9 529 18
rect 544 47 579 54
rect 544 18 554 47
rect 571 18 579 47
rect 544 9 579 18
rect 606 46 639 54
rect 606 17 614 46
rect 631 17 639 46
rect 606 9 639 17
rect 654 47 690 54
rect 654 18 665 47
rect 682 18 690 47
rect 654 9 690 18
rect 718 46 754 54
rect 718 17 726 46
rect 744 17 754 46
rect 718 9 754 17
rect 769 45 806 54
rect 769 16 779 45
rect 797 16 806 45
rect 769 9 806 16
rect 833 46 868 53
rect 833 17 841 46
rect 859 17 868 46
rect 833 9 868 17
rect 883 46 918 53
rect 883 17 892 46
rect 910 17 918 46
rect 883 9 918 17
rect 949 45 984 53
rect 949 16 957 45
rect 975 16 984 45
rect 949 9 984 16
rect 999 45 1034 53
rect 999 16 1008 45
rect 1025 16 1034 45
rect 999 9 1034 16
rect 1049 46 1084 53
rect 1049 17 1058 46
rect 1075 17 1084 46
rect 1049 9 1084 17
rect 1099 46 1134 53
rect 1099 17 1108 46
rect 1125 17 1134 46
rect 1099 9 1134 17
rect 1149 46 1187 53
rect 1149 17 1160 46
rect 1177 17 1187 46
rect 1149 9 1187 17
rect 1219 46 1253 54
rect 1219 17 1228 46
rect 1245 17 1253 46
rect 1219 9 1253 17
rect 1268 45 1303 54
rect 1268 16 1278 45
rect 1295 16 1303 45
rect 1268 9 1303 16
rect 1330 47 1365 54
rect 1330 18 1338 47
rect 1355 18 1365 47
rect 1330 9 1365 18
rect 1380 47 1415 54
rect 1380 18 1389 47
rect 1406 18 1415 47
rect 1380 9 1415 18
rect 1430 47 1465 54
rect 1430 18 1440 47
rect 1457 18 1465 47
rect 1430 9 1465 18
rect 1492 46 1525 54
rect 1492 17 1500 46
rect 1517 17 1525 46
rect 1492 9 1525 17
rect 1540 47 1576 54
rect 1540 18 1551 47
rect 1568 18 1576 47
rect 1540 9 1576 18
rect 1603 47 1639 54
rect 1603 18 1613 47
rect 1630 18 1639 47
rect 1603 9 1639 18
rect 1654 9 1691 54
rect 1706 47 1742 54
rect 1706 18 1716 47
rect 1733 18 1742 47
rect 1706 9 1742 18
rect 1779 46 1815 54
rect 1779 17 1787 46
rect 1805 17 1815 46
rect 1779 9 1815 17
rect 1830 45 1867 54
rect 1830 16 1840 45
rect 1858 16 1867 45
rect 1830 9 1867 16
<< ndiffc >>
rect -159 -133 -142 -105
rect -106 -133 -89 -105
rect -43 -138 -26 -110
rect 6 -138 23 -110
rect 72 -137 89 -109
rect 172 -138 189 -110
rect 271 -138 288 -110
rect 343 -133 360 -105
rect 392 -133 409 -105
rect 454 -133 471 -105
rect 553 -133 570 -105
rect 614 -133 631 -105
rect 664 -133 681 -105
rect 727 -133 744 -105
rect 780 -133 797 -105
rect 843 -138 860 -110
rect 892 -138 909 -110
rect 958 -137 975 -109
rect 1058 -138 1075 -110
rect 1157 -138 1174 -110
rect 1229 -133 1246 -105
rect 1278 -133 1295 -105
rect 1340 -133 1357 -105
rect 1439 -133 1456 -105
rect 1500 -133 1517 -105
rect 1550 -133 1567 -105
rect 1614 -133 1631 -105
rect 1664 -133 1681 -105
rect 1718 -133 1735 -105
rect 1788 -133 1805 -105
rect 1841 -133 1858 -105
<< pdiffc >>
rect -160 17 -142 46
rect -107 16 -89 45
rect -45 17 -27 46
rect 6 17 24 46
rect 71 16 89 45
rect 122 16 139 45
rect 172 17 189 46
rect 222 17 239 46
rect 274 17 291 46
rect 342 17 359 46
rect 392 16 409 45
rect 451 17 468 46
rect 503 18 520 47
rect 554 18 571 47
rect 614 17 631 46
rect 665 18 682 47
rect 726 17 744 46
rect 779 16 797 45
rect 841 17 859 46
rect 892 17 910 46
rect 957 16 975 45
rect 1008 16 1025 45
rect 1058 17 1075 46
rect 1108 17 1125 46
rect 1160 17 1177 46
rect 1228 17 1245 46
rect 1278 16 1295 45
rect 1338 18 1355 47
rect 1389 18 1406 47
rect 1440 18 1457 47
rect 1500 17 1517 46
rect 1551 18 1568 47
rect 1613 18 1630 47
rect 1716 18 1733 47
rect 1787 17 1805 46
rect 1840 16 1858 45
<< psubdiff >>
rect -189 -187 1892 -186
rect -189 -190 1647 -187
rect -189 -208 -122 -190
rect -105 -191 422 -190
rect -105 -208 -10 -191
rect -189 -209 -10 -208
rect 7 -209 28 -191
rect 45 -209 108 -191
rect 125 -209 151 -191
rect 168 -209 194 -191
rect 211 -209 237 -191
rect 254 -209 305 -191
rect 322 -209 387 -191
rect 404 -208 422 -191
rect 439 -191 764 -190
rect 439 -208 490 -191
rect 404 -209 490 -208
rect 507 -209 532 -191
rect 549 -209 574 -191
rect 591 -209 659 -191
rect 676 -208 764 -191
rect 781 -191 1308 -190
rect 781 -208 876 -191
rect 676 -209 876 -208
rect 893 -209 914 -191
rect 931 -209 994 -191
rect 1011 -209 1037 -191
rect 1054 -209 1080 -191
rect 1097 -209 1123 -191
rect 1140 -209 1191 -191
rect 1208 -209 1273 -191
rect 1290 -208 1308 -191
rect 1325 -191 1647 -190
rect 1325 -208 1376 -191
rect 1290 -209 1376 -208
rect 1393 -209 1418 -191
rect 1435 -209 1460 -191
rect 1477 -209 1545 -191
rect 1562 -192 1647 -191
rect 1562 -209 1579 -192
rect -189 -210 1579 -209
rect 1596 -205 1647 -192
rect 1664 -189 1892 -187
rect 1664 -191 1751 -189
rect 1664 -205 1682 -191
rect 1596 -209 1682 -205
rect 1699 -207 1751 -191
rect 1768 -207 1819 -189
rect 1836 -190 1892 -189
rect 1836 -207 1853 -190
rect 1699 -208 1853 -207
rect 1870 -208 1892 -190
rect 1699 -209 1892 -208
rect 1596 -210 1892 -209
rect -189 -215 1892 -210
<< nsubdiff >>
rect -173 122 685 125
rect -173 121 379 122
rect -173 103 -122 121
rect -105 119 24 121
rect -105 103 -12 119
rect -173 101 -12 103
rect 5 103 24 119
rect 41 120 94 121
rect 41 103 60 120
rect 5 102 60 103
rect 77 103 94 120
rect 111 103 162 121
rect 179 120 313 121
rect 179 103 200 120
rect 77 102 200 103
rect 217 119 276 120
rect 217 102 240 119
rect 5 101 240 102
rect 257 102 276 119
rect 293 103 313 120
rect 330 104 379 121
rect 396 104 417 122
rect 434 121 685 122
rect 434 120 586 121
rect 434 104 491 120
rect 330 103 491 104
rect 293 102 491 103
rect 508 102 527 120
rect 544 103 586 120
rect 603 103 642 121
rect 659 103 685 121
rect 544 102 685 103
rect 257 101 685 102
rect -173 96 685 101
rect 713 123 1875 125
rect 713 122 1723 123
rect 713 121 1265 122
rect 713 103 764 121
rect 781 119 910 121
rect 781 103 874 119
rect 713 101 874 103
rect 891 103 910 119
rect 927 120 980 121
rect 927 103 946 120
rect 891 102 946 103
rect 963 103 980 120
rect 997 103 1048 121
rect 1065 120 1199 121
rect 1065 103 1086 120
rect 963 102 1086 103
rect 1103 119 1162 120
rect 1103 102 1126 119
rect 891 101 1126 102
rect 1143 102 1162 119
rect 1179 103 1199 120
rect 1216 104 1265 121
rect 1282 104 1303 122
rect 1320 121 1654 122
rect 1320 120 1472 121
rect 1320 104 1377 120
rect 1216 103 1377 104
rect 1179 102 1377 103
rect 1394 102 1413 120
rect 1430 103 1472 120
rect 1489 103 1528 121
rect 1545 103 1569 121
rect 1586 104 1654 121
rect 1671 121 1723 122
rect 1671 104 1689 121
rect 1586 103 1689 104
rect 1706 105 1723 121
rect 1740 122 1875 123
rect 1740 121 1811 122
rect 1740 105 1757 121
rect 1706 103 1757 105
rect 1774 104 1811 121
rect 1828 104 1846 122
rect 1863 104 1875 122
rect 1774 103 1875 104
rect 1430 102 1875 103
rect 1143 101 1875 102
rect 713 96 1875 101
<< psubdiffcont >>
rect -122 -208 -105 -190
rect -10 -209 7 -191
rect 28 -209 45 -191
rect 108 -209 125 -191
rect 151 -209 168 -191
rect 194 -209 211 -191
rect 237 -209 254 -191
rect 305 -209 322 -191
rect 387 -209 404 -191
rect 422 -208 439 -190
rect 490 -209 507 -191
rect 532 -209 549 -191
rect 574 -209 591 -191
rect 659 -209 676 -191
rect 764 -208 781 -190
rect 876 -209 893 -191
rect 914 -209 931 -191
rect 994 -209 1011 -191
rect 1037 -209 1054 -191
rect 1080 -209 1097 -191
rect 1123 -209 1140 -191
rect 1191 -209 1208 -191
rect 1273 -209 1290 -191
rect 1308 -208 1325 -190
rect 1376 -209 1393 -191
rect 1418 -209 1435 -191
rect 1460 -209 1477 -191
rect 1545 -209 1562 -191
rect 1579 -210 1596 -192
rect 1647 -205 1664 -187
rect 1682 -209 1699 -191
rect 1751 -207 1768 -189
rect 1819 -207 1836 -189
rect 1853 -208 1870 -190
<< nsubdiffcont >>
rect -122 103 -105 121
rect -12 101 5 119
rect 24 103 41 121
rect 60 102 77 120
rect 94 103 111 121
rect 162 103 179 121
rect 200 102 217 120
rect 240 101 257 119
rect 276 102 293 120
rect 313 103 330 121
rect 379 104 396 122
rect 417 104 434 122
rect 491 102 508 120
rect 527 102 544 120
rect 586 103 603 121
rect 642 103 659 121
rect 764 103 781 121
rect 874 101 891 119
rect 910 103 927 121
rect 946 102 963 120
rect 980 103 997 121
rect 1048 103 1065 121
rect 1086 102 1103 120
rect 1126 101 1143 119
rect 1162 102 1179 120
rect 1199 103 1216 121
rect 1265 104 1282 122
rect 1303 104 1320 122
rect 1377 102 1394 120
rect 1413 102 1430 120
rect 1472 103 1489 121
rect 1528 103 1545 121
rect 1569 103 1586 121
rect 1654 104 1671 122
rect 1689 103 1706 121
rect 1723 105 1740 123
rect 1757 103 1774 121
rect 1811 104 1828 122
rect 1846 104 1863 122
<< poly >>
rect -132 54 -117 75
rect -18 53 -3 75
rect 98 53 113 75
rect 148 53 163 75
rect 198 53 213 75
rect 248 53 263 75
rect 367 54 382 75
rect 479 54 494 79
rect 529 54 544 79
rect 639 54 654 79
rect 754 54 769 75
rect 868 53 883 75
rect 984 53 999 75
rect 1034 53 1049 75
rect 1084 53 1099 75
rect 1134 53 1149 75
rect 1253 54 1268 75
rect 1365 54 1380 79
rect 1415 54 1430 79
rect 1525 54 1540 79
rect 1639 54 1654 79
rect 1691 54 1706 79
rect 1815 54 1830 75
rect -132 -99 -117 9
rect -18 -102 -3 9
rect 44 -61 77 -54
rect 98 -61 113 9
rect 44 -78 52 -61
rect 69 -76 113 -61
rect 69 -78 77 -76
rect 44 -85 77 -78
rect 98 -102 113 -76
rect 148 -102 163 9
rect 198 -12 213 9
rect 184 -20 213 -12
rect 184 -37 189 -20
rect 206 -37 213 -20
rect 184 -45 213 -37
rect 198 -102 213 -45
rect 248 -102 263 9
rect 313 -56 346 -49
rect 313 -73 321 -56
rect 338 -63 346 -56
rect 367 -63 382 9
rect 338 -73 382 -63
rect 313 -80 382 -73
rect 367 -97 382 -80
rect 479 -97 494 9
rect 529 -97 544 9
rect 585 -55 618 -49
rect 585 -72 593 -55
rect 610 -63 618 -55
rect 639 -63 654 9
rect 754 -10 769 9
rect 729 -15 769 -10
rect 729 -32 737 -15
rect 754 -32 769 -15
rect 729 -39 769 -32
rect 610 -72 654 -63
rect 585 -80 654 -72
rect 639 -97 654 -80
rect -132 -158 -117 -141
rect 754 -99 769 -39
rect 868 -102 883 9
rect 930 -61 963 -54
rect 984 -61 999 9
rect 930 -78 938 -61
rect 955 -76 999 -61
rect 955 -78 963 -76
rect 930 -85 963 -78
rect 984 -102 999 -76
rect 1034 -102 1049 9
rect 1084 -12 1099 9
rect 1070 -20 1099 -12
rect 1070 -37 1075 -20
rect 1092 -37 1099 -20
rect 1070 -45 1099 -37
rect 1084 -102 1099 -45
rect 1134 -15 1149 9
rect 1170 -15 1205 -10
rect 1134 -32 1178 -15
rect 1195 -32 1205 -15
rect 1134 -102 1149 -32
rect 1170 -40 1205 -32
rect 1253 -53 1268 9
rect 1365 -9 1380 9
rect 1330 -15 1380 -9
rect 1330 -32 1342 -15
rect 1359 -32 1380 -15
rect 1330 -40 1380 -32
rect 1230 -58 1268 -53
rect 1230 -75 1238 -58
rect 1255 -75 1268 -58
rect 1230 -80 1268 -75
rect 1253 -97 1268 -80
rect 1365 -97 1380 -40
rect 1415 -97 1430 9
rect 1471 -55 1504 -49
rect 1471 -72 1479 -55
rect 1496 -63 1504 -55
rect 1525 -63 1540 9
rect 1639 -42 1654 9
rect 1691 -8 1706 9
rect 1675 -16 1706 -8
rect 1675 -33 1682 -16
rect 1700 -33 1706 -16
rect 1675 -41 1706 -33
rect 1496 -72 1540 -63
rect 1471 -80 1540 -72
rect 1604 -50 1654 -42
rect 1604 -70 1612 -50
rect 1635 -70 1654 -50
rect 1604 -78 1654 -70
rect 1525 -97 1540 -80
rect 1639 -97 1654 -78
rect 1691 -97 1706 -41
rect 1815 -48 1830 9
rect 1789 -56 1830 -48
rect 1789 -73 1797 -56
rect 1815 -73 1830 -56
rect 1789 -81 1830 -73
rect -18 -160 -3 -147
rect 98 -159 113 -146
rect 148 -159 163 -146
rect 198 -159 213 -146
rect 248 -159 263 -146
rect 367 -154 382 -141
rect 479 -154 494 -141
rect 529 -154 544 -141
rect 639 -154 654 -141
rect 754 -158 769 -141
rect 1815 -99 1830 -81
rect 868 -160 883 -147
rect 984 -159 999 -146
rect 1034 -159 1049 -146
rect 1084 -159 1099 -146
rect 1134 -159 1149 -146
rect 1253 -154 1268 -141
rect 1365 -154 1380 -141
rect 1415 -154 1430 -141
rect 1525 -154 1540 -141
rect 1639 -154 1654 -141
rect 1691 -154 1706 -141
rect 1815 -158 1830 -141
<< polycont >>
rect 52 -78 69 -61
rect 189 -37 206 -20
rect 321 -73 338 -56
rect 593 -72 610 -55
rect 737 -32 754 -15
rect 938 -78 955 -61
rect 1075 -37 1092 -20
rect 1178 -32 1195 -15
rect 1342 -32 1359 -15
rect 1238 -75 1255 -58
rect 1479 -72 1496 -55
rect 1682 -33 1700 -16
rect 1612 -70 1635 -50
rect 1797 -73 1815 -56
<< locali >>
rect -191 123 1891 125
rect -191 122 1723 123
rect -191 121 122 122
rect -191 103 -161 121
rect -144 103 -122 121
rect -105 119 24 121
rect -105 103 -82 119
rect -191 101 -82 103
rect -65 101 -46 119
rect -29 101 -12 119
rect 5 103 24 119
rect 41 120 94 121
rect 41 103 60 120
rect 5 102 60 103
rect 77 103 94 120
rect 111 104 122 121
rect 139 121 343 122
rect 139 104 162 121
rect 111 103 162 104
rect 179 120 313 121
rect 179 103 200 120
rect 77 102 200 103
rect 217 119 276 120
rect 217 102 240 119
rect 5 101 240 102
rect 257 102 276 119
rect 293 103 313 120
rect 330 104 343 121
rect 360 104 379 122
rect 396 104 417 122
rect 434 121 1008 122
rect 434 120 586 121
rect 434 104 451 120
rect 330 103 451 104
rect 293 102 451 103
rect 468 102 491 120
rect 508 102 527 120
rect 544 102 552 120
rect 569 103 586 120
rect 603 120 642 121
rect 603 103 613 120
rect 569 102 613 103
rect 630 103 642 120
rect 659 103 725 121
rect 742 103 764 121
rect 781 119 910 121
rect 781 103 804 119
rect 630 102 804 103
rect 257 101 804 102
rect 821 101 840 119
rect 857 101 874 119
rect 891 103 910 119
rect 927 120 980 121
rect 927 103 946 120
rect 891 102 946 103
rect 963 103 980 120
rect 997 104 1008 121
rect 1025 121 1229 122
rect 1025 104 1048 121
rect 997 103 1048 104
rect 1065 120 1199 121
rect 1065 103 1086 120
rect 963 102 1086 103
rect 1103 119 1162 120
rect 1103 102 1126 119
rect 891 101 1126 102
rect 1143 102 1162 119
rect 1179 103 1199 120
rect 1216 104 1229 121
rect 1246 104 1265 122
rect 1282 104 1303 122
rect 1320 121 1654 122
rect 1320 120 1472 121
rect 1320 104 1337 120
rect 1216 103 1337 104
rect 1179 102 1337 103
rect 1354 102 1377 120
rect 1394 102 1413 120
rect 1430 102 1438 120
rect 1455 103 1472 120
rect 1489 120 1528 121
rect 1489 103 1499 120
rect 1455 102 1499 103
rect 1516 103 1528 120
rect 1545 103 1569 121
rect 1586 103 1616 121
rect 1633 104 1654 121
rect 1671 121 1723 122
rect 1671 104 1689 121
rect 1633 103 1689 104
rect 1706 105 1723 121
rect 1740 122 1891 123
rect 1740 121 1811 122
rect 1740 105 1757 121
rect 1706 103 1757 105
rect 1774 103 1785 121
rect 1802 104 1811 121
rect 1828 104 1846 122
rect 1863 104 1891 122
rect 1802 103 1891 104
rect 1516 102 1891 103
rect 1143 101 1891 102
rect -191 96 1891 101
rect -162 54 -143 96
rect -168 46 -134 54
rect -168 17 -160 46
rect -142 17 -134 46
rect -168 9 -134 17
rect -115 45 -80 54
rect -43 53 -26 96
rect 123 53 140 96
rect 344 54 361 96
rect 451 54 468 96
rect 554 54 571 96
rect 614 54 631 96
rect 724 54 743 96
rect -115 16 -107 45
rect -89 16 -80 45
rect -115 9 -80 16
rect -53 46 -19 53
rect -53 17 -45 46
rect -27 17 -19 46
rect -53 9 -19 17
rect -2 46 32 53
rect -2 17 6 46
rect 24 17 32 46
rect -2 9 32 17
rect 63 45 97 53
rect 63 16 71 45
rect 89 16 97 45
rect 63 9 97 16
rect 114 45 147 53
rect 114 16 122 45
rect 139 16 147 45
rect 114 9 147 16
rect 164 46 197 53
rect 164 17 172 46
rect 189 17 197 46
rect 164 9 197 17
rect 214 46 247 53
rect 214 17 222 46
rect 239 17 247 46
rect 214 9 247 17
rect 264 46 301 53
rect 264 17 274 46
rect 291 17 301 46
rect 264 9 301 17
rect 333 46 366 54
rect 333 17 342 46
rect 359 17 366 46
rect 333 9 366 17
rect 383 45 417 54
rect 383 16 392 45
rect 409 16 417 45
rect 383 9 417 16
rect 444 46 478 54
rect 444 17 451 46
rect 468 17 478 46
rect 444 9 478 17
rect 495 47 528 54
rect 495 18 503 47
rect 520 18 528 47
rect 495 9 528 18
rect 545 47 579 54
rect 545 18 554 47
rect 571 18 579 47
rect 545 9 579 18
rect 606 46 638 54
rect 606 17 614 46
rect 631 17 638 46
rect 606 9 638 17
rect 655 47 690 54
rect 655 18 665 47
rect 682 18 690 47
rect 655 9 690 18
rect 718 46 752 54
rect 718 17 726 46
rect 744 17 752 46
rect 718 9 752 17
rect 771 45 806 54
rect 843 53 860 96
rect 1009 53 1026 96
rect 1230 54 1247 96
rect 1337 54 1354 96
rect 1440 54 1457 96
rect 1500 54 1517 96
rect 1613 54 1631 96
rect 1785 54 1804 96
rect 771 16 779 45
rect 797 16 806 45
rect 771 9 806 16
rect 833 46 867 53
rect 833 17 841 46
rect 859 17 867 46
rect 833 9 867 17
rect 884 46 918 53
rect 884 17 892 46
rect 910 17 918 46
rect 884 9 918 17
rect 949 45 983 53
rect 949 16 957 45
rect 975 16 983 45
rect 949 9 983 16
rect 1000 45 1033 53
rect 1000 16 1008 45
rect 1025 16 1033 45
rect 1000 9 1033 16
rect 1050 46 1083 53
rect 1050 17 1058 46
rect 1075 17 1083 46
rect 1050 9 1083 17
rect 1100 46 1133 53
rect 1100 17 1108 46
rect 1125 17 1133 46
rect 1100 9 1133 17
rect 1150 46 1187 53
rect 1150 17 1160 46
rect 1177 17 1187 46
rect 1150 9 1187 17
rect 1219 46 1252 54
rect 1219 17 1228 46
rect 1245 17 1252 46
rect 1219 9 1252 17
rect 1269 45 1303 54
rect 1269 16 1278 45
rect 1295 16 1303 45
rect 1269 9 1303 16
rect 1330 47 1364 54
rect 1330 18 1338 47
rect 1355 18 1364 47
rect 1330 9 1364 18
rect 1381 47 1414 54
rect 1381 18 1389 47
rect 1406 18 1414 47
rect 1381 9 1414 18
rect 1431 47 1465 54
rect 1431 18 1440 47
rect 1457 18 1465 47
rect 1431 9 1465 18
rect 1492 46 1524 54
rect 1492 17 1500 46
rect 1517 17 1524 46
rect 1492 9 1524 17
rect 1541 47 1576 54
rect 1541 18 1551 47
rect 1568 18 1576 47
rect 1541 9 1576 18
rect 1603 47 1638 54
rect 1603 18 1613 47
rect 1630 18 1638 47
rect 1603 9 1638 18
rect 1707 47 1742 54
rect 1707 18 1716 47
rect 1733 18 1742 47
rect 1707 9 1742 18
rect 1779 46 1813 54
rect 1779 17 1787 46
rect 1805 17 1813 46
rect 1779 9 1813 17
rect 1832 45 1867 54
rect 1832 16 1840 45
rect 1858 16 1867 45
rect 1832 9 1867 16
rect -107 -63 -89 9
rect 7 -20 24 9
rect 184 -20 213 -12
rect 7 -37 189 -20
rect 206 -37 213 -20
rect -62 -63 -32 -57
rect -107 -80 -55 -63
rect -38 -80 -32 -63
rect -107 -99 -89 -80
rect -62 -85 -32 -80
rect -168 -105 -134 -99
rect -168 -133 -159 -105
rect -142 -133 -134 -105
rect -168 -141 -134 -133
rect -115 -105 -81 -99
rect 7 -102 24 -37
rect 184 -45 213 -37
rect 44 -61 77 -54
rect 44 -78 52 -61
rect 69 -78 77 -61
rect 230 -63 247 9
rect 395 -8 412 9
rect 387 -14 420 -8
rect 387 -31 396 -14
rect 413 -31 420 -14
rect 387 -40 420 -31
rect 313 -56 346 -49
rect 313 -63 321 -56
rect 44 -85 77 -78
rect 171 -73 321 -63
rect 338 -73 346 -56
rect 171 -80 346 -73
rect 171 -102 188 -80
rect 395 -97 412 -40
rect 502 -63 519 9
rect 665 -39 682 9
rect 729 -15 762 -10
rect 729 -32 737 -15
rect 754 -32 762 -15
rect 729 -39 762 -32
rect 585 -55 618 -49
rect 585 -63 593 -55
rect 502 -72 593 -63
rect 610 -72 618 -55
rect 502 -80 618 -72
rect 663 -53 704 -39
rect 663 -70 675 -53
rect 692 -70 704 -53
rect 663 -79 704 -70
rect 779 -63 797 9
rect 893 -20 910 9
rect 1070 -20 1099 -12
rect 893 -37 1075 -20
rect 1092 -37 1099 -20
rect 824 -63 854 -57
rect 553 -97 570 -80
rect 665 -97 682 -79
rect 779 -80 831 -63
rect 848 -80 854 -63
rect -115 -133 -106 -105
rect -89 -133 -81 -105
rect -115 -141 -81 -133
rect -53 -110 -19 -102
rect -53 -138 -43 -110
rect -26 -138 -19 -110
rect -159 -186 -142 -141
rect -53 -147 -19 -138
rect -2 -110 32 -102
rect -2 -138 6 -110
rect 23 -138 32 -110
rect -2 -147 32 -138
rect 64 -109 97 -102
rect 64 -137 72 -109
rect 89 -137 97 -109
rect 64 -146 97 -137
rect 164 -110 195 -102
rect 164 -138 172 -110
rect 189 -138 195 -110
rect 164 -146 195 -138
rect 264 -110 295 -102
rect 264 -138 271 -110
rect 288 -138 295 -110
rect 264 -146 295 -138
rect 333 -105 366 -97
rect 333 -133 343 -105
rect 360 -133 366 -105
rect 333 -141 366 -133
rect 383 -105 416 -97
rect 383 -133 392 -105
rect 409 -133 416 -105
rect 383 -141 416 -133
rect 446 -105 478 -97
rect 446 -133 454 -105
rect 471 -133 478 -105
rect 446 -141 478 -133
rect 545 -105 579 -97
rect 545 -133 553 -105
rect 570 -133 579 -105
rect 545 -141 579 -133
rect 606 -105 638 -97
rect 606 -133 614 -105
rect 631 -133 638 -105
rect 606 -141 638 -133
rect 656 -105 688 -97
rect 779 -99 797 -80
rect 824 -85 854 -80
rect 656 -133 664 -105
rect 681 -133 688 -105
rect 656 -141 688 -133
rect 718 -105 752 -99
rect 718 -133 727 -105
rect 744 -133 752 -105
rect 718 -141 752 -133
rect 771 -105 805 -99
rect 893 -102 910 -37
rect 1070 -45 1099 -37
rect 930 -61 963 -54
rect 930 -78 938 -61
rect 955 -78 963 -61
rect 1116 -63 1133 9
rect 1170 -15 1205 -10
rect 1170 -32 1178 -15
rect 1195 -32 1205 -15
rect 1170 -40 1205 -32
rect 1281 -40 1298 9
rect 1330 -15 1367 -9
rect 1330 -32 1342 -15
rect 1359 -32 1367 -15
rect 1330 -40 1367 -32
rect 1230 -58 1263 -53
rect 1230 -63 1238 -58
rect 930 -85 963 -78
rect 1057 -75 1238 -63
rect 1255 -75 1263 -58
rect 1057 -80 1263 -75
rect 1281 -57 1313 -40
rect 1057 -102 1074 -80
rect 1281 -97 1298 -57
rect 1388 -63 1405 9
rect 1551 -8 1568 9
rect 1551 -16 1706 -8
rect 1551 -25 1682 -16
rect 1471 -55 1504 -49
rect 1471 -63 1479 -55
rect 1388 -72 1479 -63
rect 1496 -72 1504 -55
rect 1388 -80 1504 -72
rect 1439 -97 1456 -80
rect 1551 -97 1568 -25
rect 1672 -33 1682 -25
rect 1700 -33 1706 -16
rect 1672 -41 1706 -33
rect 1604 -50 1643 -42
rect 1604 -70 1612 -50
rect 1635 -70 1643 -50
rect 1723 -62 1741 9
rect 1789 -56 1823 -48
rect 1789 -62 1797 -56
rect 1604 -78 1643 -70
rect 1664 -73 1797 -62
rect 1815 -73 1823 -56
rect 1664 -80 1823 -73
rect 1664 -97 1681 -80
rect 1789 -81 1823 -80
rect 1840 -63 1858 9
rect 1840 -80 1872 -63
rect 771 -133 780 -105
rect 797 -133 805 -105
rect 771 -141 805 -133
rect 833 -110 867 -102
rect 833 -138 843 -110
rect 860 -138 867 -110
rect -43 -186 -26 -147
rect 71 -186 88 -146
rect 270 -186 287 -146
rect 343 -186 360 -141
rect 454 -186 471 -141
rect 614 -186 631 -141
rect 727 -186 744 -141
rect 833 -147 867 -138
rect 884 -110 918 -102
rect 884 -138 892 -110
rect 909 -138 918 -110
rect 884 -147 918 -138
rect 950 -109 983 -102
rect 950 -137 958 -109
rect 975 -137 983 -109
rect 950 -146 983 -137
rect 1050 -110 1081 -102
rect 1050 -138 1058 -110
rect 1075 -138 1081 -110
rect 1050 -146 1081 -138
rect 1150 -110 1181 -102
rect 1150 -138 1157 -110
rect 1174 -138 1181 -110
rect 1150 -146 1181 -138
rect 1219 -105 1252 -97
rect 1219 -133 1229 -105
rect 1246 -133 1252 -105
rect 1219 -141 1252 -133
rect 1269 -105 1302 -97
rect 1269 -133 1278 -105
rect 1295 -133 1302 -105
rect 1269 -141 1302 -133
rect 1332 -105 1364 -97
rect 1332 -133 1340 -105
rect 1357 -133 1364 -105
rect 1332 -141 1364 -133
rect 1431 -105 1465 -97
rect 1431 -133 1439 -105
rect 1456 -133 1465 -105
rect 1431 -141 1465 -133
rect 1492 -105 1524 -97
rect 1492 -133 1500 -105
rect 1517 -133 1524 -105
rect 1492 -141 1524 -133
rect 1542 -105 1574 -97
rect 1542 -133 1550 -105
rect 1567 -133 1574 -105
rect 1542 -141 1574 -133
rect 1605 -105 1638 -97
rect 1605 -133 1614 -105
rect 1631 -133 1638 -105
rect 1605 -141 1638 -133
rect 1656 -105 1689 -97
rect 1656 -133 1664 -105
rect 1681 -133 1689 -105
rect 1656 -141 1689 -133
rect 1707 -105 1740 -97
rect 1840 -99 1858 -80
rect 1707 -133 1718 -105
rect 1735 -133 1740 -105
rect 1707 -141 1740 -133
rect 1779 -105 1813 -99
rect 1779 -133 1788 -105
rect 1805 -133 1813 -105
rect 1779 -141 1813 -133
rect 1832 -105 1866 -99
rect 1832 -133 1841 -105
rect 1858 -133 1866 -105
rect 1832 -141 1866 -133
rect 843 -186 860 -147
rect 957 -186 974 -146
rect 1156 -186 1173 -146
rect 1229 -186 1246 -141
rect 1340 -186 1357 -141
rect 1500 -186 1517 -141
rect 1614 -186 1631 -141
rect 1718 -186 1735 -141
rect 1788 -186 1805 -141
rect -189 -187 1892 -186
rect -189 -190 1647 -187
rect -189 -191 -122 -190
rect -189 -209 -160 -191
rect -143 -208 -122 -191
rect -105 -191 422 -190
rect -105 -208 -83 -191
rect -143 -209 -83 -208
rect -66 -209 -42 -191
rect -25 -209 -10 -191
rect 7 -209 28 -191
rect 45 -209 71 -191
rect 88 -209 108 -191
rect 125 -209 151 -191
rect 168 -209 194 -191
rect 211 -209 237 -191
rect 254 -209 269 -191
rect 286 -209 305 -191
rect 322 -209 343 -191
rect 360 -209 387 -191
rect 404 -208 422 -191
rect 439 -191 614 -190
rect 439 -208 454 -191
rect 404 -209 454 -208
rect 471 -209 490 -191
rect 507 -209 532 -191
rect 549 -209 574 -191
rect 591 -208 614 -191
rect 631 -191 764 -190
rect 631 -208 659 -191
rect 591 -209 659 -208
rect 676 -209 726 -191
rect 743 -208 764 -191
rect 781 -191 1308 -190
rect 781 -208 803 -191
rect 743 -209 803 -208
rect 820 -209 844 -191
rect 861 -209 876 -191
rect 893 -209 914 -191
rect 931 -209 957 -191
rect 974 -209 994 -191
rect 1011 -209 1037 -191
rect 1054 -209 1080 -191
rect 1097 -209 1123 -191
rect 1140 -209 1155 -191
rect 1172 -209 1191 -191
rect 1208 -209 1229 -191
rect 1246 -209 1273 -191
rect 1290 -208 1308 -191
rect 1325 -191 1500 -190
rect 1325 -208 1340 -191
rect 1290 -209 1340 -208
rect 1357 -209 1376 -191
rect 1393 -209 1418 -191
rect 1435 -209 1460 -191
rect 1477 -208 1500 -191
rect 1517 -191 1613 -190
rect 1517 -208 1545 -191
rect 1477 -209 1545 -208
rect 1562 -192 1613 -191
rect 1562 -209 1579 -192
rect -189 -210 1579 -209
rect 1596 -208 1613 -192
rect 1630 -205 1647 -190
rect 1664 -189 1892 -187
rect 1664 -191 1717 -189
rect 1664 -205 1682 -191
rect 1630 -208 1682 -205
rect 1596 -209 1682 -208
rect 1699 -207 1717 -191
rect 1734 -207 1751 -189
rect 1768 -207 1788 -189
rect 1805 -207 1819 -189
rect 1836 -190 1892 -189
rect 1836 -207 1853 -190
rect 1699 -208 1853 -207
rect 1870 -208 1892 -190
rect 1699 -209 1892 -208
rect 1596 -210 1892 -209
rect -189 -215 1892 -210
<< viali >>
rect -161 103 -144 121
rect -82 101 -65 119
rect -46 101 -29 119
rect 122 104 139 122
rect 343 104 360 122
rect 451 102 468 120
rect 552 102 569 120
rect 613 102 630 120
rect 725 103 742 121
rect 804 101 821 119
rect 840 101 857 119
rect 1008 104 1025 122
rect 1229 104 1246 122
rect 1337 102 1354 120
rect 1438 102 1455 120
rect 1499 102 1516 120
rect 1616 103 1633 121
rect 1785 103 1802 121
rect 71 16 88 45
rect 172 17 189 46
rect 274 17 291 46
rect 957 16 974 45
rect 1058 17 1075 46
rect 1160 17 1177 46
rect -55 -80 -38 -63
rect 52 -78 69 -61
rect 396 -31 413 -14
rect 737 -32 754 -15
rect 675 -70 692 -53
rect 831 -80 848 -63
rect 938 -78 955 -61
rect 1178 -32 1195 -15
rect 1342 -32 1359 -15
rect 1612 -70 1635 -50
rect -160 -209 -143 -191
rect -83 -209 -66 -191
rect -42 -209 -25 -191
rect 71 -209 88 -191
rect 269 -209 286 -191
rect 343 -209 360 -191
rect 454 -209 471 -191
rect 614 -208 631 -190
rect 726 -209 743 -191
rect 803 -209 820 -191
rect 844 -209 861 -191
rect 957 -209 974 -191
rect 1155 -209 1172 -191
rect 1229 -209 1246 -191
rect 1340 -209 1357 -191
rect 1500 -208 1517 -190
rect 1613 -208 1630 -190
rect 1717 -207 1734 -189
rect 1788 -207 1805 -189
<< metal1 >>
rect -191 122 1891 125
rect -191 121 122 122
rect -191 103 -161 121
rect -144 119 122 121
rect -144 103 -82 119
rect -191 101 -82 103
rect -65 101 -46 119
rect -29 104 122 119
rect 139 104 343 122
rect 360 121 1008 122
rect 360 120 725 121
rect 360 104 451 120
rect -29 102 451 104
rect 468 102 552 120
rect 569 102 613 120
rect 630 103 725 120
rect 742 119 1008 121
rect 742 103 804 119
rect 630 102 804 103
rect -29 101 804 102
rect 821 101 840 119
rect 857 104 1008 119
rect 1025 104 1229 122
rect 1246 121 1891 122
rect 1246 120 1616 121
rect 1246 104 1337 120
rect 857 102 1337 104
rect 1354 102 1438 120
rect 1455 102 1499 120
rect 1516 103 1616 120
rect 1633 103 1785 121
rect 1802 103 1891 121
rect 1516 102 1891 103
rect 857 101 1891 102
rect -191 96 1891 101
rect 63 45 97 53
rect 63 16 71 45
rect 88 38 97 45
rect 164 46 197 53
rect 164 38 172 46
rect 88 20 172 38
rect 88 16 97 20
rect 63 9 97 16
rect 164 17 172 20
rect 189 38 197 46
rect 264 46 301 53
rect 264 38 274 46
rect 189 20 274 38
rect 189 17 197 20
rect 164 9 197 17
rect 264 17 274 20
rect 291 17 301 46
rect 264 9 301 17
rect 949 45 983 53
rect 949 16 957 45
rect 974 38 983 45
rect 1050 46 1083 53
rect 1050 38 1058 46
rect 974 20 1058 38
rect 974 16 983 20
rect 949 9 983 16
rect 1050 17 1058 20
rect 1075 38 1083 46
rect 1150 46 1187 53
rect 1150 38 1160 46
rect 1075 20 1160 38
rect 1075 17 1083 20
rect 1050 9 1083 17
rect 1150 17 1160 20
rect 1177 17 1187 46
rect 1150 9 1187 17
rect 387 -14 420 -7
rect 387 -31 396 -14
rect 413 -15 420 -14
rect 729 -15 762 -10
rect 1170 -15 1205 -10
rect 413 -30 737 -15
rect 413 -31 420 -30
rect 387 -40 420 -31
rect 729 -32 737 -30
rect 754 -32 1178 -15
rect 1195 -18 1205 -15
rect 1330 -15 1367 -9
rect 1330 -18 1342 -15
rect 1195 -32 1342 -18
rect 1359 -32 1367 -15
rect 729 -39 762 -32
rect 1170 -40 1205 -32
rect 1330 -40 1367 -32
rect 665 -45 704 -44
rect -62 -63 -32 -57
rect 44 -61 77 -54
rect 44 -63 52 -61
rect -62 -80 -55 -63
rect -38 -78 52 -63
rect 69 -78 77 -61
rect 665 -71 672 -45
rect 698 -71 704 -45
rect 1604 -45 1643 -42
rect 665 -78 704 -71
rect 824 -63 854 -57
rect 930 -61 963 -54
rect 930 -63 938 -61
rect -38 -80 -32 -78
rect -62 -85 -32 -80
rect 44 -85 77 -78
rect 824 -80 831 -63
rect 848 -78 938 -63
rect 955 -78 963 -61
rect 1604 -72 1611 -45
rect 1638 -72 1643 -45
rect 1604 -78 1643 -72
rect 848 -80 854 -78
rect 824 -85 854 -80
rect 930 -85 963 -78
rect -189 -189 1892 -186
rect -189 -190 1717 -189
rect -189 -191 614 -190
rect -189 -209 -160 -191
rect -143 -209 -83 -191
rect -66 -209 -42 -191
rect -25 -209 71 -191
rect 88 -209 269 -191
rect 286 -209 343 -191
rect 360 -209 454 -191
rect 471 -208 614 -191
rect 631 -191 1500 -190
rect 631 -208 726 -191
rect 471 -209 726 -208
rect 743 -209 803 -191
rect 820 -209 844 -191
rect 861 -209 957 -191
rect 974 -209 1155 -191
rect 1172 -209 1229 -191
rect 1246 -209 1340 -191
rect 1357 -208 1500 -191
rect 1517 -208 1613 -190
rect 1630 -207 1717 -190
rect 1734 -207 1788 -189
rect 1805 -207 1892 -189
rect 1630 -208 1892 -207
rect 1357 -209 1892 -208
rect -189 -215 1892 -209
<< via1 >>
rect 672 -53 698 -45
rect 672 -70 675 -53
rect 675 -70 692 -53
rect 692 -70 698 -53
rect 672 -71 698 -70
rect 1611 -50 1638 -45
rect 1611 -70 1612 -50
rect 1612 -70 1635 -50
rect 1635 -70 1638 -50
rect 1611 -72 1638 -70
<< metal2 >>
rect 665 -45 704 -40
rect 665 -71 672 -45
rect 698 -57 704 -45
rect 1604 -45 1643 -42
rect 1604 -57 1611 -45
rect 698 -71 1611 -57
rect 665 -78 704 -71
rect 1604 -72 1611 -71
rect 1638 -72 1643 -45
rect 1604 -78 1643 -72
<< labels >>
flabel metal1 s -187 -211 -163 -191 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel poly s -138 -163 -114 -143 0 FreeSans 80 0 0 0 A
port 2 nsew
flabel poly s 243 -167 267 -147 0 FreeSans 80 0 0 0 A
flabel poly s -21 -167 3 -147 0 FreeSans 80 0 0 0 B
port 3 nsew
flabel poly s 144 -167 168 -147 0 FreeSans 80 0 0 0 B
flabel poly s 475 -155 498 -142 0 FreeSans 80 0 0 0 A
flabel poly s 527 -156 550 -143 0 FreeSans 80 0 0 0 B
flabel metal1 s 699 -211 723 -191 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel poly s 867 -165 886 -150 0 FreeSans 80 0 0 0 Cin
port 4 nsew
flabel poly s 1032 -161 1051 -146 0 FreeSans 80 0 0 0 Cin
flabel locali s 1303 -53 1322 -38 0 FreeSans 80 0 0 0 SUM
port 5 nsew
flabel locali s 1851 -78 1870 -63 0 FreeSans 80 0 0 0 COUT
port 6 nsew
flabel poly s 1412 -158 1435 -140 0 FreeSans 80 0 0 0 Cin
flabel metal1 s 697 100 721 120 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel metal1 s -189 100 -165 120 0 FreeSans 80 0 0 0 VDD
port 0 nsew
<< end >>
